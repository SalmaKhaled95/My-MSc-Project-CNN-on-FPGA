module TB_bla();

reg clk;
reg rst_Controller;
//reg L0START;
//wire L0FINISH;
reg [65:0] DataIn0 , DataIn1 , DataIn2 , DataIn3 ;

localparam period = 100; 
/* wire [65:0] FinalAnswer; */
wire [3:0] FinalAnswer;
//LAYER0 TheLayer(clk ,L0START, L0FINISH , DataIn0 , DataIn1 , DataIn2 , DataIn3 , DataOut0 , DataOut1 , DataOut2 , DataOut3 , DataOut4 , DataOut5 , DataOut6 , DataOut7 , DataOut8 , DataOut9 , DataOut10 , DataOut11 , DataOut12 , DataOut13 , DataOut14 , DataOut15 , DataOut16 , DataOut17 , DataOut18 , DataOut19 , DataOut20 , DataOut21 , DataOut22 , DataOut23 , DataOut24 , DataOut25 , DataOut26 , DataOut27 , DataOut28 , DataOut29 , DataOut30 , DataOut31 , DataOut32 , DataOut33 , DataOut34 , DataOut35 , DataOut36 , DataOut37 , DataOut38 , DataOut39 , DataOut40 , DataOut41 , DataOut42 , DataOut43 , DataOut44 , DataOut45 , DataOut46 , DataOut47 , DataOut48 , DataOut49 , DataOut50 , DataOut51 , DataOut52 , DataOut53 , DataOut54 , DataOut55 , DataOut56 , DataOut57 , DataOut58 , DataOut59 , DataOut60 , DataOut61 , DataOut62 , DataOut63 , DataOut64 , DataOut65 , DataOut66 , DataOut67 , DataOut68 , DataOut69 , DataOut70 , DataOut71 , DataOut72 , DataOut73 , DataOut74 , DataOut75 , DataOut76 , DataOut77 , DataOut78 , DataOut79 , DataOut80 , DataOut81 , DataOut82 , DataOut83 , DataOut84 , DataOut85 , DataOut86 , DataOut87 , DataOut88 , DataOut89 , DataOut90 , DataOut91 , DataOut92 , DataOut93 , DataOut94 , DataOut95 , DataOut96 , DataOut97 , DataOut98 , DataOut99 , DataOut100 , DataOut101 , DataOut102 , DataOut103 , DataOut104 , DataOut105 , DataOut106 , DataOut107 , DataOut108 , DataOut109 , DataOut110 , DataOut111 , DataOut112 , DataOut113 , DataOut114 , DataOut115 , DataOut116 , DataOut117 , DataOut118 , DataOut119 , DataOut120 , DataOut121 , DataOut122 , DataOut123 , DataOut124 , DataOut125 , DataOut126 , DataOut127 , DataOut128 , DataOut129 , DataOut130 , DataOut131 , DataOut132 , DataOut133 , DataOut134 , DataOut135 , DataOut136 , DataOut137 , DataOut138 , DataOut139 , DataOut140 , DataOut141 , DataOut142 , DataOut143 , DataOut144 , DataOut145 , DataOut146 , DataOut147 , DataOut148 , DataOut149 , DataOut150 , DataOut151 , DataOut152 , DataOut153 , DataOut154 , DataOut155 , DataOut156 , DataOut157 , DataOut158 , DataOut159 , DataOut160 , DataOut161 , DataOut162 , DataOut163 , DataOut164 , DataOut165 , DataOut166 , DataOut167 , DataOut168 , DataOut169 , DataOut170 , DataOut171 , DataOut172 , DataOut173 , DataOut174 , DataOut175 , DataOut176 , DataOut177 , DataOut178 , DataOut179 , DataOut180 , DataOut181 , DataOut182 , DataOut183 , DataOut184 , DataOut185 , DataOut186 , DataOut187 , DataOut188 , DataOut189 , DataOut190 , DataOut191 , DataOut192 , DataOut193 , DataOut194 , DataOut195 , DataOut196 , DataOut197 , DataOut198 , DataOut199 , DataOut200 , DataOut201 , DataOut202 , DataOut203 , DataOut204 , DataOut205 , DataOut206 , DataOut207 , DataOut208 , DataOut209 , DataOut210 , DataOut211 , DataOut212 , DataOut213 , DataOut214 , DataOut215 , DataOut216 , DataOut217 , DataOut218 , DataOut219 , DataOut220 , DataOut221 , DataOut222 , DataOut223 , DataOut224 , DataOut225 , DataOut226 , DataOut227 , DataOut228 , DataOut229 , DataOut230 , DataOut231 , DataOut232 , DataOut233 , DataOut234 , DataOut235 , DataOut236 , DataOut237 , DataOut238 , DataOut239 , DataOut240 , DataOut241 , DataOut242 , DataOut243 , DataOut244 , DataOut245 , DataOut246 , DataOut247 , DataOut248 , DataOut249 , DataOut250 , DataOut251 , DataOut252 , DataOut253 , DataOut254 , DataOut255 , DataOut256 , DataOut257 , DataOut258 , DataOut259 , DataOut260 , DataOut261 , DataOut262 , DataOut263 , DataOut264 , DataOut265 , DataOut266 , DataOut267 , DataOut268 , DataOut269 , DataOut270 , DataOut271 , DataOut272 , DataOut273 , DataOut274 , DataOut275 , DataOut276 , DataOut277 , DataOut278 , DataOut279 , DataOut280 , DataOut281 , DataOut282 , DataOut283 , DataOut284 , DataOut285 , DataOut286 , DataOut287 , DataOut288 , DataOut289 , DataOut290 , DataOut291 , DataOut292 , DataOut293 , DataOut294 , DataOut295 , DataOut296 , DataOut297 , DataOut298 , DataOut299 , DataOut300 , DataOut301 , DataOut302 , DataOut303 , DataOut304 , DataOut305 , DataOut306 , DataOut307 , DataOut308 , DataOut309 , DataOut310 , DataOut311 , DataOut312 , DataOut313 , DataOut314 , DataOut315 , DataOut316 , DataOut317 , DataOut318 , DataOut319 , DataOut320 , DataOut321 , DataOut322 , DataOut323 , DataOut324 , DataOut325 , DataOut326 , DataOut327 , DataOut328 , DataOut329 , DataOut330 , DataOut331 , DataOut332 , DataOut333 , DataOut334 , DataOut335 , DataOut336 , DataOut337 , DataOut338 , DataOut339 , DataOut340 , DataOut341 , DataOut342 , DataOut343 , DataOut344 , DataOut345 , DataOut346 , DataOut347 , DataOut348 , DataOut349 , DataOut350 , DataOut351 , DataOut352 , DataOut353 , DataOut354 , DataOut355 , DataOut356 , DataOut357 , DataOut358 , DataOut359 , DataOut360 , DataOut361 , DataOut362 , DataOut363 , DataOut364 , DataOut365 , DataOut366 , DataOut367 , DataOut368 , DataOut369 , DataOut370 , DataOut371 , DataOut372 , DataOut373 , DataOut374 , DataOut375 , DataOut376 , DataOut377 , DataOut378 , DataOut379 , DataOut380 , DataOut381 , DataOut382 , DataOut383 , DataOut384 , DataOut385 , DataOut386 , DataOut387 , DataOut388 , DataOut389 , DataOut390 , DataOut391 , DataOut392 , DataOut393 , DataOut394 , DataOut395 , DataOut396 , DataOut397 , DataOut398 , DataOut399 , DataOut400 , DataOut401 , DataOut402 , DataOut403 , DataOut404 , DataOut405 , DataOut406 , DataOut407 , DataOut408 , DataOut409 , DataOut410 , DataOut411 , DataOut412 , DataOut413 , DataOut414 , DataOut415 , DataOut416 , DataOut417 , DataOut418 , DataOut419 , DataOut420 , DataOut421 , DataOut422 , DataOut423 , DataOut424 , DataOut425 , DataOut426 , DataOut427 , DataOut428 , DataOut429 , DataOut430 , DataOut431 , DataOut432 , DataOut433 , DataOut434 , DataOut435 , DataOut436 , DataOut437 , DataOut438 , DataOut439 , DataOut440 , DataOut441 , DataOut442 , DataOut443 , DataOut444 , DataOut445 , DataOut446 , DataOut447 , DataOut448 , DataOut449 , DataOut450 , DataOut451 , DataOut452 , DataOut453 , DataOut454 , DataOut455 , DataOut456 , DataOut457 , DataOut458 , DataOut459 , DataOut460 , DataOut461 , DataOut462 , DataOut463 , DataOut464 , DataOut465 , DataOut466 , DataOut467 , DataOut468 , DataOut469 , DataOut470 , DataOut471 , DataOut472 , DataOut473 , DataOut474 , DataOut475 , DataOut476 , DataOut477 , DataOut478 , DataOut479 , DataOut480 , DataOut481 , DataOut482 , DataOut483 , DataOut484 , DataOut485 , DataOut486 , DataOut487 , DataOut488 , DataOut489 , DataOut490 , DataOut491 , DataOut492 , DataOut493 , DataOut494 , DataOut495 , DataOut496 , DataOut497 , DataOut498 , DataOut499 , DataOut500 , DataOut501 , DataOut502 , DataOut503 , DataOut504 , DataOut505 , DataOut506 , DataOut507 , DataOut508 , DataOut509 , DataOut510 , DataOut511 , DataOut512 , DataOut513 , DataOut514 , DataOut515 , DataOut516 , DataOut517 , DataOut518 , DataOut519 , DataOut520 , DataOut521 , DataOut522 , DataOut523 , DataOut524 , DataOut525 , DataOut526 , DataOut527 , DataOut528 , DataOut529 , DataOut530 , DataOut531 , DataOut532 , DataOut533 , DataOut534 , DataOut535 , DataOut536 , DataOut537 , DataOut538 , DataOut539 , DataOut540 , DataOut541 , DataOut542 , DataOut543 , DataOut544 , DataOut545 , DataOut546 , DataOut547 , DataOut548 , DataOut549 , DataOut550 , DataOut551 , DataOut552 , DataOut553 , DataOut554 , DataOut555 , DataOut556 , DataOut557 , DataOut558 , DataOut559 , DataOut560 , DataOut561 , DataOut562 , DataOut563 , DataOut564 , DataOut565 , DataOut566 , DataOut567 , DataOut568 , DataOut569 , DataOut570 , DataOut571 , DataOut572 , DataOut573 , DataOut574 , DataOut575 , DataOut576 , DataOut577 , DataOut578 , DataOut579 , DataOut580 , DataOut581 , DataOut582 , DataOut583 , DataOut584 , DataOut585 , DataOut586 , DataOut587 , DataOut588 , DataOut589 , DataOut590 , DataOut591 , DataOut592 , DataOut593 , DataOut594 , DataOut595 , DataOut596 , DataOut597 , DataOut598 , DataOut599 , DataOut600 , DataOut601 , DataOut602 , DataOut603 , DataOut604 , DataOut605 , DataOut606 , DataOut607 , DataOut608 , DataOut609 , DataOut610 , DataOut611 , DataOut612 , DataOut613 , DataOut614 , DataOut615 , DataOut616 , DataOut617 , DataOut618 , DataOut619 , DataOut620 , DataOut621 , DataOut622 , DataOut623 , DataOut624 , DataOut625 , DataOut626 , DataOut627 , DataOut628 , DataOut629 , DataOut630 , DataOut631 , DataOut632 , DataOut633 , DataOut634 , DataOut635 , DataOut636 , DataOut637 , DataOut638 , DataOut639 , DataOut640 , DataOut641 , DataOut642 , DataOut643 , DataOut644 , DataOut645 , DataOut646 , DataOut647 , DataOut648 , DataOut649 , DataOut650 , DataOut651 , DataOut652 , DataOut653 , DataOut654 , DataOut655 , DataOut656 , DataOut657 , DataOut658 , DataOut659 , DataOut660 , DataOut661 , DataOut662 , DataOut663 , DataOut664 , DataOut665 , DataOut666 , DataOut667 , DataOut668 , DataOut669 , DataOut670 , DataOut671 , DataOut672 , DataOut673 , DataOut674 , DataOut675 , DataOut676 , DataOut677 , DataOut678 , DataOut679 , DataOut680 , DataOut681 , DataOut682 , DataOut683 , DataOut684 , DataOut685 , DataOut686 , DataOut687 , DataOut688 , DataOut689 , DataOut690 , DataOut691 , DataOut692 , DataOut693 , DataOut694 , DataOut695 , DataOut696 , DataOut697 , DataOut698 , DataOut699 , DataOut700 , DataOut701 , DataOut702 , DataOut703 , DataOut704 , DataOut705 , DataOut706 , DataOut707 , DataOut708 , DataOut709 , DataOut710 , DataOut711 , DataOut712 , DataOut713 , DataOut714 , DataOut715 , DataOut716 , DataOut717 , DataOut718 , DataOut719 , DataOut720 , DataOut721 , DataOut722 , DataOut723 , DataOut724 , DataOut725 , DataOut726 , DataOut727 , DataOut728 , DataOut729 , DataOut730 , DataOut731 , DataOut732 , DataOut733 , DataOut734 , DataOut735 , DataOut736 , DataOut737 , DataOut738 , DataOut739 , DataOut740 , DataOut741 , DataOut742 , DataOut743 , DataOut744 , DataOut745 , DataOut746 , DataOut747 , DataOut748 , DataOut749 , DataOut750 , DataOut751 , DataOut752 , DataOut753 , DataOut754 , DataOut755 , DataOut756 , DataOut757 , DataOut758 , DataOut759 , DataOut760 , DataOut761 , DataOut762 , DataOut763 , DataOut764 , DataOut765 , DataOut766 , DataOut767 , DataOut768 , DataOut769 , DataOut770 , DataOut771 , DataOut772 , DataOut773 , DataOut774 , DataOut775 , DataOut776 , DataOut777 , DataOut778 , DataOut779 , DataOut780 , DataOut781 , DataOut782 , DataOut783 );
happy  otta (clk, rst_Controller,FinalAnswer,  DataIn0 , DataIn1 , DataIn2 , DataIn3);
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end

initial 
        begin
		
	    rst_Controller = 1;
		#20;
		rst_Controller = 0;
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
//repeat first input again			
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
///
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000110010000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000111110000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001100001001000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100001001000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010101100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001010010000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010011111111110000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000101010000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010101100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111010000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101011001000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101110110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100010111000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000110000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001100110011000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101100111000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001001011000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000101110000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010010000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001011010000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001001110100000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001100111111000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001011011010000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001010100110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101000111000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101110011000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010101010000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100101100000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101001010000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001100010011000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001100010011000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001000110100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000100110000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000111101000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101001000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100101011000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010011111111110000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100101110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010110010000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001010000110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111100000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101010100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001010011000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001000111100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000111101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001010100110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100011001000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010100000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101110000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000111000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000111001000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101110000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100011001000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001100111010000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000011100000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001100100110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101100000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000101000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000101100000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000111101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010010110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000110001000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000110010000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000111101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001001000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000110001000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100100011000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000111101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001001000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000110001000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010111100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101001000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000101000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000110000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101010001000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100010110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010011111111110000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000101110000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101001110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101001010000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010000100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000110101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100100001000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101110101000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000111111000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001001110000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101010100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101000010000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001001000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001001000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001000001000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001000100100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001001000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101010001000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100101011000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010101100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101110011000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101101001000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101110011000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010101100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001011100100000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101101111000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001010101100000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000100110000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000101010000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100110110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101110011000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010001100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000100000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001010011000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001100010010000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111111000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111111000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001100010010000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000110011000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000101110000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 


        end

endmodule



module LAYER0_bla (clk ,L0START, L0FINISH , DataIn0 , DataIn1 , DataIn2 , DataIn3 , DataOut0 , DataOut1 , DataOut2 , DataOut3 , DataOut4 , DataOut5 , DataOut6 , DataOut7 , DataOut8 , DataOut9 , DataOut10 , DataOut11 , DataOut12 , DataOut13 , DataOut14 , DataOut15 , DataOut16 , DataOut17 , DataOut18 , DataOut19 , DataOut20 , DataOut21 , DataOut22 , DataOut23 , DataOut24 , DataOut25 , DataOut26 , DataOut27 , DataOut28 , DataOut29 , DataOut30 , DataOut31 , DataOut32 , DataOut33 , DataOut34 , DataOut35 , DataOut36 , DataOut37 , DataOut38 , DataOut39 , DataOut40 , DataOut41 , DataOut42 , DataOut43 , DataOut44 , DataOut45 , DataOut46 , DataOut47 , DataOut48 , DataOut49 , DataOut50 , DataOut51 , DataOut52 , DataOut53 , DataOut54 , DataOut55 , DataOut56 , DataOut57 , DataOut58 , DataOut59 , DataOut60 , DataOut61 , DataOut62 , DataOut63 , DataOut64 , DataOut65 , DataOut66 , DataOut67 , DataOut68 , DataOut69 , DataOut70 , DataOut71 , DataOut72 , DataOut73 , DataOut74 , DataOut75 , DataOut76 , DataOut77 , DataOut78 , DataOut79 , DataOut80 , DataOut81 , DataOut82 , DataOut83 , DataOut84 , DataOut85 , DataOut86 , DataOut87 , DataOut88 , DataOut89 , DataOut90 , DataOut91 , DataOut92 , DataOut93 , DataOut94 , DataOut95 , DataOut96 , DataOut97 , DataOut98 , DataOut99 , DataOut100 , DataOut101 , DataOut102 , DataOut103 , DataOut104 , DataOut105 , DataOut106 , DataOut107 , DataOut108 , DataOut109 , DataOut110 , DataOut111 , DataOut112 , DataOut113 , DataOut114 , DataOut115 , DataOut116 , DataOut117 , DataOut118 , DataOut119 , DataOut120 , DataOut121 , DataOut122 , DataOut123 , DataOut124 , DataOut125 , DataOut126 , DataOut127 , DataOut128 , DataOut129 , DataOut130 , DataOut131 , DataOut132 , DataOut133 , DataOut134 , DataOut135 , DataOut136 , DataOut137 , DataOut138 , DataOut139 , DataOut140 , DataOut141 , DataOut142 , DataOut143 , DataOut144 , DataOut145 , DataOut146 , DataOut147 , DataOut148 , DataOut149 , DataOut150 , DataOut151 , DataOut152 , DataOut153 , DataOut154 , DataOut155 , DataOut156 , DataOut157 , DataOut158 , DataOut159 , DataOut160 , DataOut161 , DataOut162 , DataOut163 , DataOut164 , DataOut165 , DataOut166 , DataOut167 , DataOut168 , DataOut169 , DataOut170 , DataOut171 , DataOut172 , DataOut173 , DataOut174 , DataOut175 , DataOut176 , DataOut177 , DataOut178 , DataOut179 , DataOut180 , DataOut181 , DataOut182 , DataOut183 , DataOut184 , DataOut185 , DataOut186 , DataOut187 , DataOut188 , DataOut189 , DataOut190 , DataOut191 , DataOut192 , DataOut193 , DataOut194 , DataOut195 , DataOut196 , DataOut197 , DataOut198 , DataOut199 , DataOut200 , DataOut201 , DataOut202 , DataOut203 , DataOut204 , DataOut205 , DataOut206 , DataOut207 , DataOut208 , DataOut209 , DataOut210 , DataOut211 , DataOut212 , DataOut213 , DataOut214 , DataOut215 , DataOut216 , DataOut217 , DataOut218 , DataOut219 , DataOut220 , DataOut221 , DataOut222 , DataOut223 , DataOut224 , DataOut225 , DataOut226 , DataOut227 , DataOut228 , DataOut229 , DataOut230 , DataOut231 , DataOut232 , DataOut233 , DataOut234 , DataOut235 , DataOut236 , DataOut237 , DataOut238 , DataOut239 , DataOut240 , DataOut241 , DataOut242 , DataOut243 , DataOut244 , DataOut245 , DataOut246 , DataOut247 , DataOut248 , DataOut249 , DataOut250 , DataOut251 , DataOut252 , DataOut253 , DataOut254 , DataOut255 , DataOut256 , DataOut257 , DataOut258 , DataOut259 , DataOut260 , DataOut261 , DataOut262 , DataOut263 , DataOut264 , DataOut265 , DataOut266 , DataOut267 , DataOut268 , DataOut269 , DataOut270 , DataOut271 , DataOut272 , DataOut273 , DataOut274 , DataOut275 , DataOut276 , DataOut277 , DataOut278 , DataOut279 , DataOut280 , DataOut281 , DataOut282 , DataOut283 , DataOut284 , DataOut285 , DataOut286 , DataOut287 , DataOut288 , DataOut289 , DataOut290 , DataOut291 , DataOut292 , DataOut293 , DataOut294 , DataOut295 , DataOut296 , DataOut297 , DataOut298 , DataOut299 , DataOut300 , DataOut301 , DataOut302 , DataOut303 , DataOut304 , DataOut305 , DataOut306 , DataOut307 , DataOut308 , DataOut309 , DataOut310 , DataOut311 , DataOut312 , DataOut313 , DataOut314 , DataOut315 , DataOut316 , DataOut317 , DataOut318 , DataOut319 , DataOut320 , DataOut321 , DataOut322 , DataOut323 , DataOut324 , DataOut325 , DataOut326 , DataOut327 , DataOut328 , DataOut329 , DataOut330 , DataOut331 , DataOut332 , DataOut333 , DataOut334 , DataOut335 , DataOut336 , DataOut337 , DataOut338 , DataOut339 , DataOut340 , DataOut341 , DataOut342 , DataOut343 , DataOut344 , DataOut345 , DataOut346 , DataOut347 , DataOut348 , DataOut349 , DataOut350 , DataOut351 , DataOut352 , DataOut353 , DataOut354 , DataOut355 , DataOut356 , DataOut357 , DataOut358 , DataOut359 , DataOut360 , DataOut361 , DataOut362 , DataOut363 , DataOut364 , DataOut365 , DataOut366 , DataOut367 , DataOut368 , DataOut369 , DataOut370 , DataOut371 , DataOut372 , DataOut373 , DataOut374 , DataOut375 , DataOut376 , DataOut377 , DataOut378 , DataOut379 , DataOut380 , DataOut381 , DataOut382 , DataOut383 , DataOut384 , DataOut385 , DataOut386 , DataOut387 , DataOut388 , DataOut389 , DataOut390 , DataOut391 , DataOut392 , DataOut393 , DataOut394 , DataOut395 , DataOut396 , DataOut397 , DataOut398 , DataOut399 , DataOut400 , DataOut401 , DataOut402 , DataOut403 , DataOut404 , DataOut405 , DataOut406 , DataOut407 , DataOut408 , DataOut409 , DataOut410 , DataOut411 , DataOut412 , DataOut413 , DataOut414 , DataOut415 , DataOut416 , DataOut417 , DataOut418 , DataOut419 , DataOut420 , DataOut421 , DataOut422 , DataOut423 , DataOut424 , DataOut425 , DataOut426 , DataOut427 , DataOut428 , DataOut429 , DataOut430 , DataOut431 , DataOut432 , DataOut433 , DataOut434 , DataOut435 , DataOut436 , DataOut437 , DataOut438 , DataOut439 , DataOut440 , DataOut441 , DataOut442 , DataOut443 , DataOut444 , DataOut445 , DataOut446 , DataOut447 , DataOut448 , DataOut449 , DataOut450 , DataOut451 , DataOut452 , DataOut453 , DataOut454 , DataOut455 , DataOut456 , DataOut457 , DataOut458 , DataOut459 , DataOut460 , DataOut461 , DataOut462 , DataOut463 , DataOut464 , DataOut465 , DataOut466 , DataOut467 , DataOut468 , DataOut469 , DataOut470 , DataOut471 , DataOut472 , DataOut473 , DataOut474 , DataOut475 , DataOut476 , DataOut477 , DataOut478 , DataOut479 , DataOut480 , DataOut481 , DataOut482 , DataOut483 , DataOut484 , DataOut485 , DataOut486 , DataOut487 , DataOut488 , DataOut489 , DataOut490 , DataOut491 , DataOut492 , DataOut493 , DataOut494 , DataOut495 , DataOut496 , DataOut497 , DataOut498 , DataOut499 , DataOut500 , DataOut501 , DataOut502 , DataOut503 , DataOut504 , DataOut505 , DataOut506 , DataOut507 , DataOut508 , DataOut509 , DataOut510 , DataOut511 , DataOut512 , DataOut513 , DataOut514 , DataOut515 , DataOut516 , DataOut517 , DataOut518 , DataOut519 , DataOut520 , DataOut521 , DataOut522 , DataOut523 , DataOut524 , DataOut525 , DataOut526 , DataOut527 , DataOut528 , DataOut529 , DataOut530 , DataOut531 , DataOut532 , DataOut533 , DataOut534 , DataOut535 , DataOut536 , DataOut537 , DataOut538 , DataOut539 , DataOut540 , DataOut541 , DataOut542 , DataOut543 , DataOut544 , DataOut545 , DataOut546 , DataOut547 , DataOut548 , DataOut549 , DataOut550 , DataOut551 , DataOut552 , DataOut553 , DataOut554 , DataOut555 , DataOut556 , DataOut557 , DataOut558 , DataOut559 , DataOut560 , DataOut561 , DataOut562 , DataOut563 , DataOut564 , DataOut565 , DataOut566 , DataOut567 , DataOut568 , DataOut569 , DataOut570 , DataOut571 , DataOut572 , DataOut573 , DataOut574 , DataOut575 , DataOut576 , DataOut577 , DataOut578 , DataOut579 , DataOut580 , DataOut581 , DataOut582 , DataOut583 , DataOut584 , DataOut585 , DataOut586 , DataOut587 , DataOut588 , DataOut589 , DataOut590 , DataOut591 , DataOut592 , DataOut593 , DataOut594 , DataOut595 , DataOut596 , DataOut597 , DataOut598 , DataOut599 , DataOut600 , DataOut601 , DataOut602 , DataOut603 , DataOut604 , DataOut605 , DataOut606 , DataOut607 , DataOut608 , DataOut609 , DataOut610 , DataOut611 , DataOut612 , DataOut613 , DataOut614 , DataOut615 , DataOut616 , DataOut617 , DataOut618 , DataOut619 , DataOut620 , DataOut621 , DataOut622 , DataOut623 , DataOut624 , DataOut625 , DataOut626 , DataOut627 , DataOut628 , DataOut629 , DataOut630 , DataOut631 , DataOut632 , DataOut633 , DataOut634 , DataOut635 , DataOut636 , DataOut637 , DataOut638 , DataOut639 , DataOut640 , DataOut641 , DataOut642 , DataOut643 , DataOut644 , DataOut645 , DataOut646 , DataOut647 , DataOut648 , DataOut649 , DataOut650 , DataOut651 , DataOut652 , DataOut653 , DataOut654 , DataOut655 , DataOut656 , DataOut657 , DataOut658 , DataOut659 , DataOut660 , DataOut661 , DataOut662 , DataOut663 , DataOut664 , DataOut665 , DataOut666 , DataOut667 , DataOut668 , DataOut669 , DataOut670 , DataOut671 , DataOut672 , DataOut673 , DataOut674 , DataOut675 , DataOut676 , DataOut677 , DataOut678 , DataOut679 , DataOut680 , DataOut681 , DataOut682 , DataOut683 , DataOut684 , DataOut685 , DataOut686 , DataOut687 , DataOut688 , DataOut689 , DataOut690 , DataOut691 , DataOut692 , DataOut693 , DataOut694 , DataOut695 , DataOut696 , DataOut697 , DataOut698 , DataOut699 , DataOut700 , DataOut701 , DataOut702 , DataOut703 , DataOut704 , DataOut705 , DataOut706 , DataOut707 , DataOut708 , DataOut709 , DataOut710 , DataOut711 , DataOut712 , DataOut713 , DataOut714 , DataOut715 , DataOut716 , DataOut717 , DataOut718 , DataOut719 , DataOut720 , DataOut721 , DataOut722 , DataOut723 , DataOut724 , DataOut725 , DataOut726 , DataOut727 , DataOut728 , DataOut729 , DataOut730 , DataOut731 , DataOut732 , DataOut733 , DataOut734 , DataOut735 , DataOut736 , DataOut737 , DataOut738 , DataOut739 , DataOut740 , DataOut741 , DataOut742 , DataOut743 , DataOut744 , DataOut745 , DataOut746 , DataOut747 , DataOut748 , DataOut749 , DataOut750 , DataOut751 , DataOut752 , DataOut753 , DataOut754 , DataOut755 , DataOut756 , DataOut757 , DataOut758 , DataOut759 , DataOut760 , DataOut761 , DataOut762 , DataOut763 , DataOut764 , DataOut765 , DataOut766 , DataOut767 , DataOut768 , DataOut769 , DataOut770 , DataOut771 , DataOut772 , DataOut773 , DataOut774 , DataOut775 , DataOut776 , DataOut777 , DataOut778 , DataOut779 , DataOut780 , DataOut781 , DataOut782 , DataOut783 );

input clk;
output reg [65:0] DataOut0 , DataOut1 , DataOut2 , DataOut3 , DataOut4 , DataOut5 , DataOut6 , DataOut7 , DataOut8 , DataOut9 , DataOut10 , DataOut11 , DataOut12 , DataOut13 , DataOut14 , DataOut15 , DataOut16 , DataOut17 , DataOut18 , DataOut19 , DataOut20 , DataOut21 , DataOut22 , DataOut23 , DataOut24 , DataOut25 , DataOut26 , DataOut27 , DataOut28 , DataOut29 , DataOut30 , DataOut31 , DataOut32 , DataOut33 , DataOut34 , DataOut35 , DataOut36 , DataOut37 , DataOut38 , DataOut39 , DataOut40 , DataOut41 , DataOut42 , DataOut43 , DataOut44 , DataOut45 , DataOut46 , DataOut47 , DataOut48 , DataOut49 , DataOut50 , DataOut51 , DataOut52 , DataOut53 , DataOut54 , DataOut55 , DataOut56 , DataOut57 , DataOut58 , DataOut59 , DataOut60 , DataOut61 , DataOut62 , DataOut63 , DataOut64 , DataOut65 , DataOut66 , DataOut67 , DataOut68 , DataOut69 , DataOut70 , DataOut71 , DataOut72 , DataOut73 , DataOut74 , DataOut75 , DataOut76 , DataOut77 , DataOut78 , DataOut79 , DataOut80 , DataOut81 , DataOut82 , DataOut83 , DataOut84 , DataOut85 , DataOut86 , DataOut87 , DataOut88 , DataOut89 , DataOut90 , DataOut91 , DataOut92 , DataOut93 , DataOut94 , DataOut95 , DataOut96 , DataOut97 , DataOut98 , DataOut99 , DataOut100 , DataOut101 , DataOut102 , DataOut103 , DataOut104 , DataOut105 , DataOut106 , DataOut107 , DataOut108 , DataOut109 , DataOut110 , DataOut111 , DataOut112 , DataOut113 , DataOut114 , DataOut115 , DataOut116 , DataOut117 , DataOut118 , DataOut119 , DataOut120 , DataOut121 , DataOut122 , DataOut123 , DataOut124 , DataOut125 , DataOut126 , DataOut127 , DataOut128 , DataOut129 , DataOut130 , DataOut131 , DataOut132 , DataOut133 , DataOut134 , DataOut135 , DataOut136 , DataOut137 , DataOut138 , DataOut139 , DataOut140 , DataOut141 , DataOut142 , DataOut143 , DataOut144 , DataOut145 , DataOut146 , DataOut147 , DataOut148 , DataOut149 , DataOut150 , DataOut151 , DataOut152 , DataOut153 , DataOut154 , DataOut155 , DataOut156 , DataOut157 , DataOut158 , DataOut159 , DataOut160 , DataOut161 , DataOut162 , DataOut163 , DataOut164 , DataOut165 , DataOut166 , DataOut167 , DataOut168 , DataOut169 , DataOut170 , DataOut171 , DataOut172 , DataOut173 , DataOut174 , DataOut175 , DataOut176 , DataOut177 , DataOut178 , DataOut179 , DataOut180 , DataOut181 , DataOut182 , DataOut183 , DataOut184 , DataOut185 , DataOut186 , DataOut187 , DataOut188 , DataOut189 , DataOut190 , DataOut191 , DataOut192 , DataOut193 , DataOut194 , DataOut195 , DataOut196 , DataOut197 , DataOut198 , DataOut199 , DataOut200 , DataOut201 , DataOut202 , DataOut203 , DataOut204 , DataOut205 , DataOut206 , DataOut207 , DataOut208 , DataOut209 , DataOut210 , DataOut211 , DataOut212 , DataOut213 , DataOut214 , DataOut215 , DataOut216 , DataOut217 , DataOut218 , DataOut219 , DataOut220 , DataOut221 , DataOut222 , DataOut223 , DataOut224 , DataOut225 , DataOut226 , DataOut227 , DataOut228 , DataOut229 , DataOut230 , DataOut231 , DataOut232 , DataOut233 , DataOut234 , DataOut235 , DataOut236 , DataOut237 , DataOut238 , DataOut239 , DataOut240 , DataOut241 , DataOut242 , DataOut243 , DataOut244 , DataOut245 , DataOut246 , DataOut247 , DataOut248 , DataOut249 , DataOut250 , DataOut251 , DataOut252 , DataOut253 , DataOut254 , DataOut255 , DataOut256 , DataOut257 , DataOut258 , DataOut259 , DataOut260 , DataOut261 , DataOut262 , DataOut263 , DataOut264 , DataOut265 , DataOut266 , DataOut267 , DataOut268 , DataOut269 , DataOut270 , DataOut271 , DataOut272 , DataOut273 , DataOut274 , DataOut275 , DataOut276 , DataOut277 , DataOut278 , DataOut279 , DataOut280 , DataOut281 , DataOut282 , DataOut283 , DataOut284 , DataOut285 , DataOut286 , DataOut287 , DataOut288 , DataOut289 , DataOut290 , DataOut291 , DataOut292 , DataOut293 , DataOut294 , DataOut295 , DataOut296 , DataOut297 , DataOut298 , DataOut299 , DataOut300 , DataOut301 , DataOut302 , DataOut303 , DataOut304 , DataOut305 , DataOut306 , DataOut307 , DataOut308 , DataOut309 , DataOut310 , DataOut311 , DataOut312 , DataOut313 , DataOut314 , DataOut315 , DataOut316 , DataOut317 , DataOut318 , DataOut319 , DataOut320 , DataOut321 , DataOut322 , DataOut323 , DataOut324 , DataOut325 , DataOut326 , DataOut327 , DataOut328 , DataOut329 , DataOut330 , DataOut331 , DataOut332 , DataOut333 , DataOut334 , DataOut335 , DataOut336 , DataOut337 , DataOut338 , DataOut339 , DataOut340 , DataOut341 , DataOut342 , DataOut343 , DataOut344 , DataOut345 , DataOut346 , DataOut347 , DataOut348 , DataOut349 , DataOut350 , DataOut351 , DataOut352 , DataOut353 , DataOut354 , DataOut355 , DataOut356 , DataOut357 , DataOut358 , DataOut359 , DataOut360 , DataOut361 , DataOut362 , DataOut363 , DataOut364 , DataOut365 , DataOut366 , DataOut367 , DataOut368 , DataOut369 , DataOut370 , DataOut371 , DataOut372 , DataOut373 , DataOut374 , DataOut375 , DataOut376 , DataOut377 , DataOut378 , DataOut379 , DataOut380 , DataOut381 , DataOut382 , DataOut383 , DataOut384 , DataOut385 , DataOut386 , DataOut387 , DataOut388 , DataOut389 , DataOut390 , DataOut391 , DataOut392 , DataOut393 , DataOut394 , DataOut395 , DataOut396 , DataOut397 , DataOut398 , DataOut399 , DataOut400 , DataOut401 , DataOut402 , DataOut403 , DataOut404 , DataOut405 , DataOut406 , DataOut407 , DataOut408 , DataOut409 , DataOut410 , DataOut411 , DataOut412 , DataOut413 , DataOut414 , DataOut415 , DataOut416 , DataOut417 , DataOut418 , DataOut419 , DataOut420 , DataOut421 , DataOut422 , DataOut423 , DataOut424 , DataOut425 , DataOut426 , DataOut427 , DataOut428 , DataOut429 , DataOut430 , DataOut431 , DataOut432 , DataOut433 , DataOut434 , DataOut435 , DataOut436 , DataOut437 , DataOut438 , DataOut439 , DataOut440 , DataOut441 , DataOut442 , DataOut443 , DataOut444 , DataOut445 , DataOut446 , DataOut447 , DataOut448 , DataOut449 , DataOut450 , DataOut451 , DataOut452 , DataOut453 , DataOut454 , DataOut455 , DataOut456 , DataOut457 , DataOut458 , DataOut459 , DataOut460 , DataOut461 , DataOut462 , DataOut463 , DataOut464 , DataOut465 , DataOut466 , DataOut467 , DataOut468 , DataOut469 , DataOut470 , DataOut471 , DataOut472 , DataOut473 , DataOut474 , DataOut475 , DataOut476 , DataOut477 , DataOut478 , DataOut479 , DataOut480 , DataOut481 , DataOut482 , DataOut483 , DataOut484 , DataOut485 , DataOut486 , DataOut487 , DataOut488 , DataOut489 , DataOut490 , DataOut491 , DataOut492 , DataOut493 , DataOut494 , DataOut495 , DataOut496 , DataOut497 , DataOut498 , DataOut499 , DataOut500 , DataOut501 , DataOut502 , DataOut503 , DataOut504 , DataOut505 , DataOut506 , DataOut507 , DataOut508 , DataOut509 , DataOut510 , DataOut511 , DataOut512 , DataOut513 , DataOut514 , DataOut515 , DataOut516 , DataOut517 , DataOut518 , DataOut519 , DataOut520 , DataOut521 , DataOut522 , DataOut523 , DataOut524 , DataOut525 , DataOut526 , DataOut527 , DataOut528 , DataOut529 , DataOut530 , DataOut531 , DataOut532 , DataOut533 , DataOut534 , DataOut535 , DataOut536 , DataOut537 , DataOut538 , DataOut539 , DataOut540 , DataOut541 , DataOut542 , DataOut543 , DataOut544 , DataOut545 , DataOut546 , DataOut547 , DataOut548 , DataOut549 , DataOut550 , DataOut551 , DataOut552 , DataOut553 , DataOut554 , DataOut555 , DataOut556 , DataOut557 , DataOut558 , DataOut559 , DataOut560 , DataOut561 , DataOut562 , DataOut563 , DataOut564 , DataOut565 , DataOut566 , DataOut567 , DataOut568 , DataOut569 , DataOut570 , DataOut571 , DataOut572 , DataOut573 , DataOut574 , DataOut575 , DataOut576 , DataOut577 , DataOut578 , DataOut579 , DataOut580 , DataOut581 , DataOut582 , DataOut583 , DataOut584 , DataOut585 , DataOut586 , DataOut587 , DataOut588 , DataOut589 , DataOut590 , DataOut591 , DataOut592 , DataOut593 , DataOut594 , DataOut595 , DataOut596 , DataOut597 , DataOut598 , DataOut599 , DataOut600 , DataOut601 , DataOut602 , DataOut603 , DataOut604 , DataOut605 , DataOut606 , DataOut607 , DataOut608 , DataOut609 , DataOut610 , DataOut611 , DataOut612 , DataOut613 , DataOut614 , DataOut615 , DataOut616 , DataOut617 , DataOut618 , DataOut619 , DataOut620 , DataOut621 , DataOut622 , DataOut623 , DataOut624 , DataOut625 , DataOut626 , DataOut627 , DataOut628 , DataOut629 , DataOut630 , DataOut631 , DataOut632 , DataOut633 , DataOut634 , DataOut635 , DataOut636 , DataOut637 , DataOut638 , DataOut639 , DataOut640 , DataOut641 , DataOut642 , DataOut643 , DataOut644 , DataOut645 , DataOut646 , DataOut647 , DataOut648 , DataOut649 , DataOut650 , DataOut651 , DataOut652 , DataOut653 , DataOut654 , DataOut655 , DataOut656 , DataOut657 , DataOut658 , DataOut659 , DataOut660 , DataOut661 , DataOut662 , DataOut663 , DataOut664 , DataOut665 , DataOut666 , DataOut667 , DataOut668 , DataOut669 , DataOut670 , DataOut671 , DataOut672 , DataOut673 , DataOut674 , DataOut675 , DataOut676 , DataOut677 , DataOut678 , DataOut679 , DataOut680 , DataOut681 , DataOut682 , DataOut683 , DataOut684 , DataOut685 , DataOut686 , DataOut687 , DataOut688 , DataOut689 , DataOut690 , DataOut691 , DataOut692 , DataOut693 , DataOut694 , DataOut695 , DataOut696 , DataOut697 , DataOut698 , DataOut699 , DataOut700 , DataOut701 , DataOut702 , DataOut703 , DataOut704 , DataOut705 , DataOut706 , DataOut707 , DataOut708 , DataOut709 , DataOut710 , DataOut711 , DataOut712 , DataOut713 , DataOut714 , DataOut715 , DataOut716 , DataOut717 , DataOut718 , DataOut719 , DataOut720 , DataOut721 , DataOut722 , DataOut723 , DataOut724 , DataOut725 , DataOut726 , DataOut727 , DataOut728 , DataOut729 , DataOut730 , DataOut731 , DataOut732 , DataOut733 , DataOut734 , DataOut735 , DataOut736 , DataOut737 , DataOut738 , DataOut739 , DataOut740 , DataOut741 , DataOut742 , DataOut743 , DataOut744 , DataOut745 , DataOut746 , DataOut747 , DataOut748 , DataOut749 , DataOut750 , DataOut751 , DataOut752 , DataOut753 , DataOut754 , DataOut755 , DataOut756 , DataOut757 , DataOut758 , DataOut759 , DataOut760 , DataOut761 , DataOut762 , DataOut763 , DataOut764 , DataOut765 , DataOut766 , DataOut767 , DataOut768 , DataOut769 , DataOut770 , DataOut771 , DataOut772 , DataOut773 , DataOut774 , DataOut775 , DataOut776 , DataOut777 , DataOut778 , DataOut779 , DataOut780 , DataOut781 , DataOut782 , DataOut783  ;
input L0START;
output reg L0FINISH;
input wire [65:0] DataIn0 , DataIn1 , DataIn2 , DataIn3 ;
wire [7:0] counter; 
wire dump; 
COUNTER_LAYER_256_cycles TheCounter (clk, counter, L0START,dump);
//counter 196 cycles : 8 bits
always @(posedge clk) 
begin 

//$monitor("counter = %b, L0START = %b, L0FINISH = %b , DataIn0= %b", counter , L0START, L0FINISH, DataIn0);

if (L0START)
begin
//$display("one");

case(counter)
0  : begin DataOut0  <=  DataIn0; DataOut1  <=  DataIn1; DataOut2  <=  DataIn2; DataOut3  <=  DataIn3; end //$display("two"); 
1  : begin DataOut4  <=  DataIn0; DataOut5  <=  DataIn1; DataOut6  <=  DataIn2; DataOut7  <=  DataIn3; end //$display("three");
2  : begin DataOut8  <=  DataIn0; DataOut9  <=  DataIn1; DataOut10  <=  DataIn2; DataOut11  <=  DataIn3; end
3  : begin DataOut12  <=  DataIn0; DataOut13  <=  DataIn1; DataOut14  <=  DataIn2; DataOut15  <=  DataIn3; end
4  : begin DataOut16  <=  DataIn0; DataOut17  <=  DataIn1; DataOut18  <=  DataIn2; DataOut19  <=  DataIn3; end
5  : begin DataOut20  <=  DataIn0; DataOut21  <=  DataIn1; DataOut22  <=  DataIn2; DataOut23  <=  DataIn3; end
6  : begin DataOut24  <=  DataIn0; DataOut25  <=  DataIn1; DataOut26  <=  DataIn2; DataOut27  <=  DataIn3; end
7  : begin DataOut28  <=  DataIn0; DataOut29  <=  DataIn1; DataOut30  <=  DataIn2; DataOut31  <=  DataIn3; end
8  : begin DataOut32  <=  DataIn0; DataOut33  <=  DataIn1; DataOut34  <=  DataIn2; DataOut35  <=  DataIn3; end
9  : begin DataOut36  <=  DataIn0; DataOut37  <=  DataIn1; DataOut38  <=  DataIn2; DataOut39  <=  DataIn3; end
10  : begin DataOut40  <=  DataIn0; DataOut41  <=  DataIn1; DataOut42  <=  DataIn2; DataOut43  <=  DataIn3; end
11  : begin DataOut44  <=  DataIn0; DataOut45  <=  DataIn1; DataOut46  <=  DataIn2; DataOut47  <=  DataIn3; end
12  : begin DataOut48  <=  DataIn0; DataOut49  <=  DataIn1; DataOut50  <=  DataIn2; DataOut51  <=  DataIn3; end
13  : begin DataOut52  <=  DataIn0; DataOut53  <=  DataIn1; DataOut54  <=  DataIn2; DataOut55  <=  DataIn3; end
14  : begin DataOut56  <=  DataIn0; DataOut57  <=  DataIn1; DataOut58  <=  DataIn2; DataOut59  <=  DataIn3; end
15  : begin DataOut60  <=  DataIn0; DataOut61  <=  DataIn1; DataOut62  <=  DataIn2; DataOut63  <=  DataIn3; end
16  : begin DataOut64  <=  DataIn0; DataOut65  <=  DataIn1; DataOut66  <=  DataIn2; DataOut67  <=  DataIn3; end
17  : begin DataOut68  <=  DataIn0; DataOut69  <=  DataIn1; DataOut70  <=  DataIn2; DataOut71  <=  DataIn3; end
18  : begin DataOut72  <=  DataIn0; DataOut73  <=  DataIn1; DataOut74  <=  DataIn2; DataOut75  <=  DataIn3; end
19  : begin DataOut76  <=  DataIn0; DataOut77  <=  DataIn1; DataOut78  <=  DataIn2; DataOut79  <=  DataIn3; end
20  : begin DataOut80  <=  DataIn0; DataOut81  <=  DataIn1; DataOut82  <=  DataIn2; DataOut83  <=  DataIn3; end
21  : begin DataOut84  <=  DataIn0; DataOut85  <=  DataIn1; DataOut86  <=  DataIn2; DataOut87  <=  DataIn3; end
22  : begin DataOut88  <=  DataIn0; DataOut89  <=  DataIn1; DataOut90  <=  DataIn2; DataOut91  <=  DataIn3; end
23  : begin DataOut92  <=  DataIn0; DataOut93  <=  DataIn1; DataOut94  <=  DataIn2; DataOut95  <=  DataIn3; end
24  : begin DataOut96  <=  DataIn0; DataOut97  <=  DataIn1; DataOut98  <=  DataIn2; DataOut99  <=  DataIn3; end
25  : begin DataOut100  <=  DataIn0; DataOut101  <=  DataIn1; DataOut102  <=  DataIn2; DataOut103  <=  DataIn3; end
26  : begin DataOut104  <=  DataIn0; DataOut105  <=  DataIn1; DataOut106  <=  DataIn2; DataOut107  <=  DataIn3; end
27  : begin DataOut108  <=  DataIn0; DataOut109  <=  DataIn1; DataOut110  <=  DataIn2; DataOut111  <=  DataIn3; end
28  : begin DataOut112  <=  DataIn0; DataOut113  <=  DataIn1; DataOut114  <=  DataIn2; DataOut115  <=  DataIn3; end
29  : begin DataOut116  <=  DataIn0; DataOut117  <=  DataIn1; DataOut118  <=  DataIn2; DataOut119  <=  DataIn3; end
30  : begin DataOut120  <=  DataIn0; DataOut121  <=  DataIn1; DataOut122  <=  DataIn2; DataOut123  <=  DataIn3; end
31  : begin DataOut124  <=  DataIn0; DataOut125  <=  DataIn1; DataOut126  <=  DataIn2; DataOut127  <=  DataIn3; end
32  : begin DataOut128  <=  DataIn0; DataOut129  <=  DataIn1; DataOut130  <=  DataIn2; DataOut131  <=  DataIn3; end
33  : begin DataOut132  <=  DataIn0; DataOut133  <=  DataIn1; DataOut134  <=  DataIn2; DataOut135  <=  DataIn3; end
34  : begin DataOut136  <=  DataIn0; DataOut137  <=  DataIn1; DataOut138  <=  DataIn2; DataOut139  <=  DataIn3; end
35  : begin DataOut140  <=  DataIn0; DataOut141  <=  DataIn1; DataOut142  <=  DataIn2; DataOut143  <=  DataIn3; end
36  : begin DataOut144  <=  DataIn0; DataOut145  <=  DataIn1; DataOut146  <=  DataIn2; DataOut147  <=  DataIn3; end
37  : begin DataOut148  <=  DataIn0; DataOut149  <=  DataIn1; DataOut150  <=  DataIn2; DataOut151  <=  DataIn3; end
38  : begin DataOut152  <=  DataIn0; DataOut153  <=  DataIn1; DataOut154  <=  DataIn2; DataOut155  <=  DataIn3; end
39  : begin DataOut156  <=  DataIn0; DataOut157  <=  DataIn1; DataOut158  <=  DataIn2; DataOut159  <=  DataIn3; end
40  : begin DataOut160  <=  DataIn0; DataOut161  <=  DataIn1; DataOut162  <=  DataIn2; DataOut163  <=  DataIn3; end
41  : begin DataOut164  <=  DataIn0; DataOut165  <=  DataIn1; DataOut166  <=  DataIn2; DataOut167  <=  DataIn3; end
42  : begin DataOut168  <=  DataIn0; DataOut169  <=  DataIn1; DataOut170  <=  DataIn2; DataOut171  <=  DataIn3; end
43  : begin DataOut172  <=  DataIn0; DataOut173  <=  DataIn1; DataOut174  <=  DataIn2; DataOut175  <=  DataIn3; end
44  : begin DataOut176  <=  DataIn0; DataOut177  <=  DataIn1; DataOut178  <=  DataIn2; DataOut179  <=  DataIn3; end
45  : begin DataOut180  <=  DataIn0; DataOut181  <=  DataIn1; DataOut182  <=  DataIn2; DataOut183  <=  DataIn3; end
46  : begin DataOut184  <=  DataIn0; DataOut185  <=  DataIn1; DataOut186  <=  DataIn2; DataOut187  <=  DataIn3; end
47  : begin DataOut188  <=  DataIn0; DataOut189  <=  DataIn1; DataOut190  <=  DataIn2; DataOut191  <=  DataIn3; end
48  : begin DataOut192  <=  DataIn0; DataOut193  <=  DataIn1; DataOut194  <=  DataIn2; DataOut195  <=  DataIn3; end
49  : begin DataOut196  <=  DataIn0; DataOut197  <=  DataIn1; DataOut198  <=  DataIn2; DataOut199  <=  DataIn3; end
50  : begin DataOut200  <=  DataIn0; DataOut201  <=  DataIn1; DataOut202  <=  DataIn2; DataOut203  <=  DataIn3; end
51  : begin DataOut204  <=  DataIn0; DataOut205  <=  DataIn1; DataOut206  <=  DataIn2; DataOut207  <=  DataIn3; end
52  : begin DataOut208  <=  DataIn0; DataOut209  <=  DataIn1; DataOut210  <=  DataIn2; DataOut211  <=  DataIn3; end
53  : begin DataOut212  <=  DataIn0; DataOut213  <=  DataIn1; DataOut214  <=  DataIn2; DataOut215  <=  DataIn3; end
54  : begin DataOut216  <=  DataIn0; DataOut217  <=  DataIn1; DataOut218  <=  DataIn2; DataOut219  <=  DataIn3; end
55  : begin DataOut220  <=  DataIn0; DataOut221  <=  DataIn1; DataOut222  <=  DataIn2; DataOut223  <=  DataIn3; end
56  : begin DataOut224  <=  DataIn0; DataOut225  <=  DataIn1; DataOut226  <=  DataIn2; DataOut227  <=  DataIn3; end
57  : begin DataOut228  <=  DataIn0; DataOut229  <=  DataIn1; DataOut230  <=  DataIn2; DataOut231  <=  DataIn3; end
58  : begin DataOut232  <=  DataIn0; DataOut233  <=  DataIn1; DataOut234  <=  DataIn2; DataOut235  <=  DataIn3; end
59  : begin DataOut236  <=  DataIn0; DataOut237  <=  DataIn1; DataOut238  <=  DataIn2; DataOut239  <=  DataIn3; end
60  : begin DataOut240  <=  DataIn0; DataOut241  <=  DataIn1; DataOut242  <=  DataIn2; DataOut243  <=  DataIn3; end
61  : begin DataOut244  <=  DataIn0; DataOut245  <=  DataIn1; DataOut246  <=  DataIn2; DataOut247  <=  DataIn3; end
62  : begin DataOut248  <=  DataIn0; DataOut249  <=  DataIn1; DataOut250  <=  DataIn2; DataOut251  <=  DataIn3; end
63  : begin DataOut252  <=  DataIn0; DataOut253  <=  DataIn1; DataOut254  <=  DataIn2; DataOut255  <=  DataIn3; end
64  : begin DataOut256  <=  DataIn0; DataOut257  <=  DataIn1; DataOut258  <=  DataIn2; DataOut259  <=  DataIn3; end
65  : begin DataOut260  <=  DataIn0; DataOut261  <=  DataIn1; DataOut262  <=  DataIn2; DataOut263  <=  DataIn3; end
66  : begin DataOut264  <=  DataIn0; DataOut265  <=  DataIn1; DataOut266  <=  DataIn2; DataOut267  <=  DataIn3; end
67  : begin DataOut268  <=  DataIn0; DataOut269  <=  DataIn1; DataOut270  <=  DataIn2; DataOut271  <=  DataIn3; end
68  : begin DataOut272  <=  DataIn0; DataOut273  <=  DataIn1; DataOut274  <=  DataIn2; DataOut275  <=  DataIn3; end
69  : begin DataOut276  <=  DataIn0; DataOut277  <=  DataIn1; DataOut278  <=  DataIn2; DataOut279  <=  DataIn3; end
70  : begin DataOut280  <=  DataIn0; DataOut281  <=  DataIn1; DataOut282  <=  DataIn2; DataOut283  <=  DataIn3; end
71  : begin DataOut284  <=  DataIn0; DataOut285  <=  DataIn1; DataOut286  <=  DataIn2; DataOut287  <=  DataIn3; end
72  : begin DataOut288  <=  DataIn0; DataOut289  <=  DataIn1; DataOut290  <=  DataIn2; DataOut291  <=  DataIn3; end
73  : begin DataOut292  <=  DataIn0; DataOut293  <=  DataIn1; DataOut294  <=  DataIn2; DataOut295  <=  DataIn3; end
74  : begin DataOut296  <=  DataIn0; DataOut297  <=  DataIn1; DataOut298  <=  DataIn2; DataOut299  <=  DataIn3; end
75  : begin DataOut300  <=  DataIn0; DataOut301  <=  DataIn1; DataOut302  <=  DataIn2; DataOut303  <=  DataIn3; end
76  : begin DataOut304  <=  DataIn0; DataOut305  <=  DataIn1; DataOut306  <=  DataIn2; DataOut307  <=  DataIn3; end
77  : begin DataOut308  <=  DataIn0; DataOut309  <=  DataIn1; DataOut310  <=  DataIn2; DataOut311  <=  DataIn3; end
78  : begin DataOut312  <=  DataIn0; DataOut313  <=  DataIn1; DataOut314  <=  DataIn2; DataOut315  <=  DataIn3; end
79  : begin DataOut316  <=  DataIn0; DataOut317  <=  DataIn1; DataOut318  <=  DataIn2; DataOut319  <=  DataIn3; end
80  : begin DataOut320  <=  DataIn0; DataOut321  <=  DataIn1; DataOut322  <=  DataIn2; DataOut323  <=  DataIn3; end
81  : begin DataOut324  <=  DataIn0; DataOut325  <=  DataIn1; DataOut326  <=  DataIn2; DataOut327  <=  DataIn3; end
82  : begin DataOut328  <=  DataIn0; DataOut329  <=  DataIn1; DataOut330  <=  DataIn2; DataOut331  <=  DataIn3; end
83  : begin DataOut332  <=  DataIn0; DataOut333  <=  DataIn1; DataOut334  <=  DataIn2; DataOut335  <=  DataIn3; end
84  : begin DataOut336  <=  DataIn0; DataOut337  <=  DataIn1; DataOut338  <=  DataIn2; DataOut339  <=  DataIn3; end
85  : begin DataOut340  <=  DataIn0; DataOut341  <=  DataIn1; DataOut342  <=  DataIn2; DataOut343  <=  DataIn3; end
86  : begin DataOut344  <=  DataIn0; DataOut345  <=  DataIn1; DataOut346  <=  DataIn2; DataOut347  <=  DataIn3; end
87  : begin DataOut348  <=  DataIn0; DataOut349  <=  DataIn1; DataOut350  <=  DataIn2; DataOut351  <=  DataIn3; end
88  : begin DataOut352  <=  DataIn0; DataOut353  <=  DataIn1; DataOut354  <=  DataIn2; DataOut355  <=  DataIn3; end
89  : begin DataOut356  <=  DataIn0; DataOut357  <=  DataIn1; DataOut358  <=  DataIn2; DataOut359  <=  DataIn3; end
90  : begin DataOut360  <=  DataIn0; DataOut361  <=  DataIn1; DataOut362  <=  DataIn2; DataOut363  <=  DataIn3; end
91  : begin DataOut364  <=  DataIn0; DataOut365  <=  DataIn1; DataOut366  <=  DataIn2; DataOut367  <=  DataIn3; end
92  : begin DataOut368  <=  DataIn0; DataOut369  <=  DataIn1; DataOut370  <=  DataIn2; DataOut371  <=  DataIn3; end
93  : begin DataOut372  <=  DataIn0; DataOut373  <=  DataIn1; DataOut374  <=  DataIn2; DataOut375  <=  DataIn3; end
94  : begin DataOut376  <=  DataIn0; DataOut377  <=  DataIn1; DataOut378  <=  DataIn2; DataOut379  <=  DataIn3; end
95  : begin DataOut380  <=  DataIn0; DataOut381  <=  DataIn1; DataOut382  <=  DataIn2; DataOut383  <=  DataIn3; end
96  : begin DataOut384  <=  DataIn0; DataOut385  <=  DataIn1; DataOut386  <=  DataIn2; DataOut387  <=  DataIn3; end
97  : begin DataOut388  <=  DataIn0; DataOut389  <=  DataIn1; DataOut390  <=  DataIn2; DataOut391  <=  DataIn3; end
98  : begin DataOut392  <=  DataIn0; DataOut393  <=  DataIn1; DataOut394  <=  DataIn2; DataOut395  <=  DataIn3; end
99  : begin DataOut396  <=  DataIn0; DataOut397  <=  DataIn1; DataOut398  <=  DataIn2; DataOut399  <=  DataIn3; end
100  : begin DataOut400  <=  DataIn0; DataOut401  <=  DataIn1; DataOut402  <=  DataIn2; DataOut403  <=  DataIn3; end
101  : begin DataOut404  <=  DataIn0; DataOut405  <=  DataIn1; DataOut406  <=  DataIn2; DataOut407  <=  DataIn3; end
102  : begin DataOut408  <=  DataIn0; DataOut409  <=  DataIn1; DataOut410  <=  DataIn2; DataOut411  <=  DataIn3; end
103  : begin DataOut412  <=  DataIn0; DataOut413  <=  DataIn1; DataOut414  <=  DataIn2; DataOut415  <=  DataIn3; end
104  : begin DataOut416  <=  DataIn0; DataOut417  <=  DataIn1; DataOut418  <=  DataIn2; DataOut419  <=  DataIn3; end
105  : begin DataOut420  <=  DataIn0; DataOut421  <=  DataIn1; DataOut422  <=  DataIn2; DataOut423  <=  DataIn3; end
106  : begin DataOut424  <=  DataIn0; DataOut425  <=  DataIn1; DataOut426  <=  DataIn2; DataOut427  <=  DataIn3; end
107  : begin DataOut428  <=  DataIn0; DataOut429  <=  DataIn1; DataOut430  <=  DataIn2; DataOut431  <=  DataIn3; end
108  : begin DataOut432  <=  DataIn0; DataOut433  <=  DataIn1; DataOut434  <=  DataIn2; DataOut435  <=  DataIn3; end
109  : begin DataOut436  <=  DataIn0; DataOut437  <=  DataIn1; DataOut438  <=  DataIn2; DataOut439  <=  DataIn3; end
110  : begin DataOut440  <=  DataIn0; DataOut441  <=  DataIn1; DataOut442  <=  DataIn2; DataOut443  <=  DataIn3; end
111  : begin DataOut444  <=  DataIn0; DataOut445  <=  DataIn1; DataOut446  <=  DataIn2; DataOut447  <=  DataIn3; end
112  : begin DataOut448  <=  DataIn0; DataOut449  <=  DataIn1; DataOut450  <=  DataIn2; DataOut451  <=  DataIn3; end
113  : begin DataOut452  <=  DataIn0; DataOut453  <=  DataIn1; DataOut454  <=  DataIn2; DataOut455  <=  DataIn3; end
114  : begin DataOut456  <=  DataIn0; DataOut457  <=  DataIn1; DataOut458  <=  DataIn2; DataOut459  <=  DataIn3; end
115  : begin DataOut460  <=  DataIn0; DataOut461  <=  DataIn1; DataOut462  <=  DataIn2; DataOut463  <=  DataIn3; end
116  : begin DataOut464  <=  DataIn0; DataOut465  <=  DataIn1; DataOut466  <=  DataIn2; DataOut467  <=  DataIn3; end
117  : begin DataOut468  <=  DataIn0; DataOut469  <=  DataIn1; DataOut470  <=  DataIn2; DataOut471  <=  DataIn3; end
118  : begin DataOut472  <=  DataIn0; DataOut473  <=  DataIn1; DataOut474  <=  DataIn2; DataOut475  <=  DataIn3; end
119  : begin DataOut476  <=  DataIn0; DataOut477  <=  DataIn1; DataOut478  <=  DataIn2; DataOut479  <=  DataIn3; end
120  : begin DataOut480  <=  DataIn0; DataOut481  <=  DataIn1; DataOut482  <=  DataIn2; DataOut483  <=  DataIn3; end
121  : begin DataOut484  <=  DataIn0; DataOut485  <=  DataIn1; DataOut486  <=  DataIn2; DataOut487  <=  DataIn3; end
122  : begin DataOut488  <=  DataIn0; DataOut489  <=  DataIn1; DataOut490  <=  DataIn2; DataOut491  <=  DataIn3; end
123  : begin DataOut492  <=  DataIn0; DataOut493  <=  DataIn1; DataOut494  <=  DataIn2; DataOut495  <=  DataIn3; end
124  : begin DataOut496  <=  DataIn0; DataOut497  <=  DataIn1; DataOut498  <=  DataIn2; DataOut499  <=  DataIn3; end
125  : begin DataOut500  <=  DataIn0; DataOut501  <=  DataIn1; DataOut502  <=  DataIn2; DataOut503  <=  DataIn3; end
126  : begin DataOut504  <=  DataIn0; DataOut505  <=  DataIn1; DataOut506  <=  DataIn2; DataOut507  <=  DataIn3; end
127  : begin DataOut508  <=  DataIn0; DataOut509  <=  DataIn1; DataOut510  <=  DataIn2; DataOut511  <=  DataIn3; end
128  : begin DataOut512  <=  DataIn0; DataOut513  <=  DataIn1; DataOut514  <=  DataIn2; DataOut515  <=  DataIn3; end
129  : begin DataOut516  <=  DataIn0; DataOut517  <=  DataIn1; DataOut518  <=  DataIn2; DataOut519  <=  DataIn3; end
130  : begin DataOut520  <=  DataIn0; DataOut521  <=  DataIn1; DataOut522  <=  DataIn2; DataOut523  <=  DataIn3; end
131  : begin DataOut524  <=  DataIn0; DataOut525  <=  DataIn1; DataOut526  <=  DataIn2; DataOut527  <=  DataIn3; end
132  : begin DataOut528  <=  DataIn0; DataOut529  <=  DataIn1; DataOut530  <=  DataIn2; DataOut531  <=  DataIn3; end
133  : begin DataOut532  <=  DataIn0; DataOut533  <=  DataIn1; DataOut534  <=  DataIn2; DataOut535  <=  DataIn3; end
134  : begin DataOut536  <=  DataIn0; DataOut537  <=  DataIn1; DataOut538  <=  DataIn2; DataOut539  <=  DataIn3; end
135  : begin DataOut540  <=  DataIn0; DataOut541  <=  DataIn1; DataOut542  <=  DataIn2; DataOut543  <=  DataIn3; end
136  : begin DataOut544  <=  DataIn0; DataOut545  <=  DataIn1; DataOut546  <=  DataIn2; DataOut547  <=  DataIn3; end
137  : begin DataOut548  <=  DataIn0; DataOut549  <=  DataIn1; DataOut550  <=  DataIn2; DataOut551  <=  DataIn3; end
138  : begin DataOut552  <=  DataIn0; DataOut553  <=  DataIn1; DataOut554  <=  DataIn2; DataOut555  <=  DataIn3; end
139  : begin DataOut556  <=  DataIn0; DataOut557  <=  DataIn1; DataOut558  <=  DataIn2; DataOut559  <=  DataIn3; end
140  : begin DataOut560  <=  DataIn0; DataOut561  <=  DataIn1; DataOut562  <=  DataIn2; DataOut563  <=  DataIn3; end
141  : begin DataOut564  <=  DataIn0; DataOut565  <=  DataIn1; DataOut566  <=  DataIn2; DataOut567  <=  DataIn3; end
142  : begin DataOut568  <=  DataIn0; DataOut569  <=  DataIn1; DataOut570  <=  DataIn2; DataOut571  <=  DataIn3; end
143  : begin DataOut572  <=  DataIn0; DataOut573  <=  DataIn1; DataOut574  <=  DataIn2; DataOut575  <=  DataIn3; end
144  : begin DataOut576  <=  DataIn0; DataOut577  <=  DataIn1; DataOut578  <=  DataIn2; DataOut579  <=  DataIn3; end
145  : begin DataOut580  <=  DataIn0; DataOut581  <=  DataIn1; DataOut582  <=  DataIn2; DataOut583  <=  DataIn3; end
146  : begin DataOut584  <=  DataIn0; DataOut585  <=  DataIn1; DataOut586  <=  DataIn2; DataOut587  <=  DataIn3; end
147  : begin DataOut588  <=  DataIn0; DataOut589  <=  DataIn1; DataOut590  <=  DataIn2; DataOut591  <=  DataIn3; end
148  : begin DataOut592  <=  DataIn0; DataOut593  <=  DataIn1; DataOut594  <=  DataIn2; DataOut595  <=  DataIn3; end
149  : begin DataOut596  <=  DataIn0; DataOut597  <=  DataIn1; DataOut598  <=  DataIn2; DataOut599  <=  DataIn3; end
150  : begin DataOut600  <=  DataIn0; DataOut601  <=  DataIn1; DataOut602  <=  DataIn2; DataOut603  <=  DataIn3; end
151  : begin DataOut604  <=  DataIn0; DataOut605  <=  DataIn1; DataOut606  <=  DataIn2; DataOut607  <=  DataIn3; end
152  : begin DataOut608  <=  DataIn0; DataOut609  <=  DataIn1; DataOut610  <=  DataIn2; DataOut611  <=  DataIn3; end
153  : begin DataOut612  <=  DataIn0; DataOut613  <=  DataIn1; DataOut614  <=  DataIn2; DataOut615  <=  DataIn3; end
154  : begin DataOut616  <=  DataIn0; DataOut617  <=  DataIn1; DataOut618  <=  DataIn2; DataOut619  <=  DataIn3; end
155  : begin DataOut620  <=  DataIn0; DataOut621  <=  DataIn1; DataOut622  <=  DataIn2; DataOut623  <=  DataIn3; end
156  : begin DataOut624  <=  DataIn0; DataOut625  <=  DataIn1; DataOut626  <=  DataIn2; DataOut627  <=  DataIn3; end
157  : begin DataOut628  <=  DataIn0; DataOut629  <=  DataIn1; DataOut630  <=  DataIn2; DataOut631  <=  DataIn3; end
158  : begin DataOut632  <=  DataIn0; DataOut633  <=  DataIn1; DataOut634  <=  DataIn2; DataOut635  <=  DataIn3; end
159  : begin DataOut636  <=  DataIn0; DataOut637  <=  DataIn1; DataOut638  <=  DataIn2; DataOut639  <=  DataIn3; end
160  : begin DataOut640  <=  DataIn0; DataOut641  <=  DataIn1; DataOut642  <=  DataIn2; DataOut643  <=  DataIn3; end
161  : begin DataOut644  <=  DataIn0; DataOut645  <=  DataIn1; DataOut646  <=  DataIn2; DataOut647  <=  DataIn3; end
162  : begin DataOut648  <=  DataIn0; DataOut649  <=  DataIn1; DataOut650  <=  DataIn2; DataOut651  <=  DataIn3; end
163  : begin DataOut652  <=  DataIn0; DataOut653  <=  DataIn1; DataOut654  <=  DataIn2; DataOut655  <=  DataIn3; end
164  : begin DataOut656  <=  DataIn0; DataOut657  <=  DataIn1; DataOut658  <=  DataIn2; DataOut659  <=  DataIn3; end
165  : begin DataOut660  <=  DataIn0; DataOut661  <=  DataIn1; DataOut662  <=  DataIn2; DataOut663  <=  DataIn3; end
166  : begin DataOut664  <=  DataIn0; DataOut665  <=  DataIn1; DataOut666  <=  DataIn2; DataOut667  <=  DataIn3; end
167  : begin DataOut668  <=  DataIn0; DataOut669  <=  DataIn1; DataOut670  <=  DataIn2; DataOut671  <=  DataIn3; end
168  : begin DataOut672  <=  DataIn0; DataOut673  <=  DataIn1; DataOut674  <=  DataIn2; DataOut675  <=  DataIn3; end
169  : begin DataOut676  <=  DataIn0; DataOut677  <=  DataIn1; DataOut678  <=  DataIn2; DataOut679  <=  DataIn3; end
170  : begin DataOut680  <=  DataIn0; DataOut681  <=  DataIn1; DataOut682  <=  DataIn2; DataOut683  <=  DataIn3; end
171  : begin DataOut684  <=  DataIn0; DataOut685  <=  DataIn1; DataOut686  <=  DataIn2; DataOut687  <=  DataIn3; end
172  : begin DataOut688  <=  DataIn0; DataOut689  <=  DataIn1; DataOut690  <=  DataIn2; DataOut691  <=  DataIn3; end
173  : begin DataOut692  <=  DataIn0; DataOut693  <=  DataIn1; DataOut694  <=  DataIn2; DataOut695  <=  DataIn3; end
174  : begin DataOut696  <=  DataIn0; DataOut697  <=  DataIn1; DataOut698  <=  DataIn2; DataOut699  <=  DataIn3; end
175  : begin DataOut700  <=  DataIn0; DataOut701  <=  DataIn1; DataOut702  <=  DataIn2; DataOut703  <=  DataIn3; end
176  : begin DataOut704  <=  DataIn0; DataOut705  <=  DataIn1; DataOut706  <=  DataIn2; DataOut707  <=  DataIn3; end
177  : begin DataOut708  <=  DataIn0; DataOut709  <=  DataIn1; DataOut710  <=  DataIn2; DataOut711  <=  DataIn3; end
178  : begin DataOut712  <=  DataIn0; DataOut713  <=  DataIn1; DataOut714  <=  DataIn2; DataOut715  <=  DataIn3; end
179  : begin DataOut716  <=  DataIn0; DataOut717  <=  DataIn1; DataOut718  <=  DataIn2; DataOut719  <=  DataIn3; end
180  : begin DataOut720  <=  DataIn0; DataOut721  <=  DataIn1; DataOut722  <=  DataIn2; DataOut723  <=  DataIn3; end
181  : begin DataOut724  <=  DataIn0; DataOut725  <=  DataIn1; DataOut726  <=  DataIn2; DataOut727  <=  DataIn3; end
182  : begin DataOut728  <=  DataIn0; DataOut729  <=  DataIn1; DataOut730  <=  DataIn2; DataOut731  <=  DataIn3; end
183  : begin DataOut732  <=  DataIn0; DataOut733  <=  DataIn1; DataOut734  <=  DataIn2; DataOut735  <=  DataIn3; end
184  : begin DataOut736  <=  DataIn0; DataOut737  <=  DataIn1; DataOut738  <=  DataIn2; DataOut739  <=  DataIn3; end
185  : begin DataOut740  <=  DataIn0; DataOut741  <=  DataIn1; DataOut742  <=  DataIn2; DataOut743  <=  DataIn3; end
186  : begin DataOut744  <=  DataIn0; DataOut745  <=  DataIn1; DataOut746  <=  DataIn2; DataOut747  <=  DataIn3; end
187  : begin DataOut748  <=  DataIn0; DataOut749  <=  DataIn1; DataOut750  <=  DataIn2; DataOut751  <=  DataIn3; end
188  : begin DataOut752  <=  DataIn0; DataOut753  <=  DataIn1; DataOut754  <=  DataIn2; DataOut755  <=  DataIn3; end
189  : begin DataOut756  <=  DataIn0; DataOut757  <=  DataIn1; DataOut758  <=  DataIn2; DataOut759  <=  DataIn3; end
190  : begin DataOut760  <=  DataIn0; DataOut761  <=  DataIn1; DataOut762  <=  DataIn2; DataOut763  <=  DataIn3; end
191  : begin DataOut764  <=  DataIn0; DataOut765  <=  DataIn1; DataOut766  <=  DataIn2; DataOut767  <=  DataIn3; end
192  : begin DataOut768  <=  DataIn0; DataOut769  <=  DataIn1; DataOut770  <=  DataIn2; DataOut771  <=  DataIn3; end
193  : begin DataOut772  <=  DataIn0; DataOut773  <=  DataIn1; DataOut774  <=  DataIn2; DataOut775  <=  DataIn3; end
194  : begin DataOut776  <=  DataIn0; DataOut777  <=  DataIn1; DataOut778  <=  DataIn2; DataOut779  <=  DataIn3; end
195  : begin DataOut780  <=  DataIn0; DataOut781  <=  DataIn1; DataOut782  <=  DataIn2; DataOut783  <=  DataIn3; end
196  : begin L0FINISH<= 1; end //$display("four");
default: begin L0FINISH<= 1; end //$display("five");


endcase
end
 //$display("six"); 
end

endmodule


