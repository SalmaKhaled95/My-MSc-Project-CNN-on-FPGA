module MERGEHOPE_L1_L2 (clk, MAX1LayerFinish, Conv1LayerStart, DataOut0 , DataOut1 , DataOut2 , DataOut3 , DataOut4 , DataOut5 , DataOut6 , DataOut7 , DataOut8 , DataOut9 , DataOut10 , DataOut11 , DataOut12 , DataOut13 , DataOut14 , DataOut15 , DataOut16 , DataOut17 , DataOut18 , DataOut19 , DataOut20 , DataOut21 , DataOut22 , DataOut23 , DataOut24 , DataOut25 , DataOut26 , DataOut27 , DataOut28 , DataOut29 , DataOut30 , DataOut31 , DataOut32 , DataOut33 , DataOut34 , DataOut35 , DataOut36 , DataOut37 , DataOut38 , DataOut39 , DataOut40 , DataOut41 , DataOut42 , DataOut43 , DataOut44 , DataOut45 , DataOut46 , DataOut47 , DataOut48 , DataOut49 , DataOut50 , DataOut51 , DataOut52 , DataOut53 , DataOut54 , DataOut55 , DataOut56 , DataOut57 , DataOut58 , DataOut59 , DataOut60 , DataOut61 , DataOut62 , DataOut63 , DataOut64 , DataOut65 , DataOut66 , DataOut67 , DataOut68 , DataOut69 , DataOut70 , DataOut71 , DataOut72 , DataOut73 , DataOut74 , DataOut75 , DataOut76 , DataOut77 , DataOut78 , DataOut79 , DataOut80 , DataOut81 , DataOut82 , DataOut83 , DataOut84 , DataOut85 , DataOut86 , DataOut87 , DataOut88 , DataOut89 , DataOut90 , DataOut91 , DataOut92 , DataOut93 , DataOut94 , DataOut95 , DataOut96 , DataOut97 , DataOut98 , DataOut99 , DataOut100 , DataOut101 , DataOut102 , DataOut103 , DataOut104 , DataOut105 , DataOut106 , DataOut107 , DataOut108 , DataOut109 , DataOut110 , DataOut111 , DataOut112 , DataOut113 , DataOut114 , DataOut115 , DataOut116 , DataOut117 , DataOut118 , DataOut119 , DataOut120 , DataOut121 , DataOut122 , DataOut123 , DataOut124 , DataOut125 , DataOut126 , DataOut127 , DataOut128 , DataOut129 , DataOut130 , DataOut131 , DataOut132 , DataOut133 , DataOut134 , DataOut135 , DataOut136 , DataOut137 , DataOut138 , DataOut139 , DataOut140 , DataOut141 , DataOut142 , DataOut143 , DataOut144 , DataOut145 , DataOut146 , DataOut147 , DataOut148 , DataOut149 , DataOut150 , DataOut151 , DataOut152 , DataOut153 , DataOut154 , DataOut155 , DataOut156 , DataOut157 , DataOut158 , DataOut159 , DataOut160 , DataOut161 , DataOut162 , DataOut163 , DataOut164 , DataOut165 , DataOut166 , DataOut167 , DataOut168 , DataOut169 , DataOut170 , DataOut171 , DataOut172 , DataOut173 , DataOut174 , DataOut175 , DataOut176 , DataOut177 , DataOut178 , DataOut179 , DataOut180 , DataOut181 , DataOut182 , DataOut183 , DataOut184 , DataOut185 , DataOut186 , DataOut187 , DataOut188 , DataOut189 , DataOut190 , DataOut191 , DataOut192 , DataOut193 , DataOut194 , DataOut195 , DataOut196 , DataOut197 , DataOut198 , DataOut199 , DataOut200 , DataOut201 , DataOut202 , DataOut203 , DataOut204 , DataOut205 , DataOut206 , DataOut207 , DataOut208 , DataOut209 , DataOut210 , DataOut211 , DataOut212 , DataOut213 , DataOut214 , DataOut215 , DataOut216 , DataOut217 , DataOut218 , DataOut219 , DataOut220 , DataOut221 , DataOut222 , DataOut223 , DataOut224 , DataOut225 , DataOut226 , DataOut227 , DataOut228 , DataOut229 , DataOut230 , DataOut231 , DataOut232 , DataOut233 , DataOut234 , DataOut235 , DataOut236 , DataOut237 , DataOut238 , DataOut239 , DataOut240 , DataOut241 , DataOut242 , DataOut243 , DataOut244 , DataOut245 , DataOut246 , DataOut247 , DataOut248 , DataOut249 , DataOut250 , DataOut251 , DataOut252 , DataOut253 , DataOut254 , DataOut255 , DataOut256 , DataOut257 , DataOut258 , DataOut259 , DataOut260 , DataOut261 , DataOut262 , DataOut263 , DataOut264 , DataOut265 , DataOut266 , DataOut267 , DataOut268 , DataOut269 , DataOut270 , DataOut271 , DataOut272 , DataOut273 , DataOut274 , DataOut275 , DataOut276 , DataOut277 , DataOut278 , DataOut279 , DataOut280 , DataOut281 , DataOut282 , DataOut283 , DataOut284 , DataOut285 , DataOut286 , DataOut287 , DataOut288 , DataOut289 , DataOut290 , DataOut291 , DataOut292 , DataOut293 , DataOut294 , DataOut295 , DataOut296 , DataOut297 , DataOut298 , DataOut299 , DataOut300 , DataOut301 , DataOut302 , DataOut303 , DataOut304 , DataOut305 , DataOut306 , DataOut307 , DataOut308 , DataOut309 , DataOut310 , DataOut311 , DataOut312 , DataOut313 , DataOut314 , DataOut315 , DataOut316 , DataOut317 , DataOut318 , DataOut319 , DataOut320 , DataOut321 , DataOut322 , DataOut323 , DataOut324 , DataOut325 , DataOut326 , DataOut327 , DataOut328 , DataOut329 , DataOut330 , DataOut331 , DataOut332 , DataOut333 , DataOut334 , DataOut335 , DataOut336 , DataOut337 , DataOut338 , DataOut339 , DataOut340 , DataOut341 , DataOut342 , DataOut343 , DataOut344 , DataOut345 , DataOut346 , DataOut347 , DataOut348 , DataOut349 , DataOut350 , DataOut351 , DataOut352 , DataOut353 , DataOut354 , DataOut355 , DataOut356 , DataOut357 , DataOut358 , DataOut359 , DataOut360 , DataOut361 , DataOut362 , DataOut363 , DataOut364 , DataOut365 , DataOut366 , DataOut367 , DataOut368 , DataOut369 , DataOut370 , DataOut371 , DataOut372 , DataOut373 , DataOut374 , DataOut375 , DataOut376 , DataOut377 , DataOut378 , DataOut379 , DataOut380 , DataOut381 , DataOut382 , DataOut383 , DataOut384 , DataOut385 , DataOut386 , DataOut387 , DataOut388 , DataOut389 , DataOut390 , DataOut391 , DataOut392 , DataOut393 , DataOut394 , DataOut395 , DataOut396 , DataOut397 , DataOut398 , DataOut399 , DataOut400 , DataOut401 , DataOut402 , DataOut403 , DataOut404 , DataOut405 , DataOut406 , DataOut407 , DataOut408 , DataOut409 , DataOut410 , DataOut411 , DataOut412 , DataOut413 , DataOut414 , DataOut415 , DataOut416 , DataOut417 , DataOut418 , DataOut419 , DataOut420 , DataOut421 , DataOut422 , DataOut423 , DataOut424 , DataOut425 , DataOut426 , DataOut427 , DataOut428 , DataOut429 , DataOut430 , DataOut431 , DataOut432 , DataOut433 , DataOut434 , DataOut435 , DataOut436 , DataOut437 , DataOut438 , DataOut439 , DataOut440 , DataOut441 , DataOut442 , DataOut443 , DataOut444 , DataOut445 , DataOut446 , DataOut447 , DataOut448 , DataOut449 , DataOut450 , DataOut451 , DataOut452 , DataOut453 , DataOut454 , DataOut455 , DataOut456 , DataOut457 , DataOut458 , DataOut459 , DataOut460 , DataOut461 , DataOut462 , DataOut463 , DataOut464 , DataOut465 , DataOut466 , DataOut467 , DataOut468 , DataOut469 , DataOut470 , DataOut471 , DataOut472 , DataOut473 , DataOut474 , DataOut475 , DataOut476 , DataOut477 , DataOut478 , DataOut479 , DataOut480 , DataOut481 , DataOut482 , DataOut483 , DataOut484 , DataOut485 , DataOut486 , DataOut487 , DataOut488 , DataOut489 , DataOut490 , DataOut491 , DataOut492 , DataOut493 , DataOut494 , DataOut495 , DataOut496 , DataOut497 , DataOut498 , DataOut499 , DataOut500 , DataOut501 , DataOut502 , DataOut503 , DataOut504 , DataOut505 , DataOut506 , DataOut507 , DataOut508 , DataOut509 , DataOut510 , DataOut511 , DataOut512 , DataOut513 , DataOut514 , DataOut515 , DataOut516 , DataOut517 , DataOut518 , DataOut519 , DataOut520 , DataOut521 , DataOut522 , DataOut523 , DataOut524 , DataOut525 , DataOut526 , DataOut527 , DataOut528 , DataOut529 , DataOut530 , DataOut531 , DataOut532 , DataOut533 , DataOut534 , DataOut535 , DataOut536 , DataOut537 , DataOut538 , DataOut539 , DataOut540 , DataOut541 , DataOut542 , DataOut543 , DataOut544 , DataOut545 , DataOut546 , DataOut547 , DataOut548 , DataOut549 , DataOut550 , DataOut551 , DataOut552 , DataOut553 , DataOut554 , DataOut555 , DataOut556 , DataOut557 , DataOut558 , DataOut559 , DataOut560 , DataOut561 , DataOut562 , DataOut563 , DataOut564 , DataOut565 , DataOut566 , DataOut567 , DataOut568 , DataOut569 , DataOut570 , DataOut571 , DataOut572 , DataOut573 , DataOut574 , DataOut575 , DataOut576 , DataOut577 , DataOut578 , DataOut579 , DataOut580 , DataOut581 , DataOut582 , DataOut583 , DataOut584 , DataOut585 , DataOut586 , DataOut587 , DataOut588 , DataOut589 , DataOut590 , DataOut591 , DataOut592 , DataOut593 , DataOut594 , DataOut595 , DataOut596 , DataOut597 , DataOut598 , DataOut599 , DataOut600 , DataOut601 , DataOut602 , DataOut603 , DataOut604 , DataOut605 , DataOut606 , DataOut607 , DataOut608 , DataOut609 , DataOut610 , DataOut611 , DataOut612 , DataOut613 , DataOut614 , DataOut615 , DataOut616 , DataOut617 , DataOut618 , DataOut619 , DataOut620 , DataOut621 , DataOut622 , DataOut623 , DataOut624 , DataOut625 , DataOut626 , DataOut627 , DataOut628 , DataOut629 , DataOut630 , DataOut631 , DataOut632 , DataOut633 , DataOut634 , DataOut635 , DataOut636 , DataOut637 , DataOut638 , DataOut639 , DataOut640 , DataOut641 , DataOut642 , DataOut643 , DataOut644 , DataOut645 , DataOut646 , DataOut647 , DataOut648 , DataOut649 , DataOut650 , DataOut651 , DataOut652 , DataOut653 , DataOut654 , DataOut655 , DataOut656 , DataOut657 , DataOut658 , DataOut659 , DataOut660 , DataOut661 , DataOut662 , DataOut663 , DataOut664 , DataOut665 , DataOut666 , DataOut667 , DataOut668 , DataOut669 , DataOut670 , DataOut671 , DataOut672 , DataOut673 , DataOut674 , DataOut675 , DataOut676 , DataOut677 , DataOut678 , DataOut679 , DataOut680 , DataOut681 , DataOut682 , DataOut683 , DataOut684 , DataOut685 , DataOut686 , DataOut687 , DataOut688 , DataOut689 , DataOut690 , DataOut691 , DataOut692 , DataOut693 , DataOut694 , DataOut695 , DataOut696 , DataOut697 , DataOut698 , DataOut699 , DataOut700 , DataOut701 , DataOut702 , DataOut703 , DataOut704 , DataOut705 , DataOut706 , DataOut707 , DataOut708 , DataOut709 , DataOut710 , DataOut711 , DataOut712 , DataOut713 , DataOut714 , DataOut715 , DataOut716 , DataOut717 , DataOut718 , DataOut719 , DataOut720 , DataOut721 , DataOut722 , DataOut723 , DataOut724 , DataOut725 , DataOut726 , DataOut727 , DataOut728 , DataOut729 , DataOut730 , DataOut731 , DataOut732 , DataOut733 , DataOut734 , DataOut735 , DataOut736 , DataOut737 , DataOut738 , DataOut739 , DataOut740 , DataOut741 , DataOut742 , DataOut743 , DataOut744 , DataOut745 , DataOut746 , DataOut747 , DataOut748 , DataOut749 , DataOut750 , DataOut751 , DataOut752 , DataOut753 , DataOut754 , DataOut755 , DataOut756 , DataOut757 , DataOut758 , DataOut759 , DataOut760 , DataOut761 , DataOut762 , DataOut763 , DataOut764 , DataOut765 , DataOut766 , DataOut767 , DataOut768 , DataOut769 , DataOut770 , DataOut771 , DataOut772 , DataOut773 , DataOut774 , DataOut775 , DataOut776 , DataOut777 , DataOut778 , DataOut779 , DataOut780 , DataOut781 , DataOut782 , DataOut783 
,REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143 
);


input clk;
input wire [65:0] DataOut0 , DataOut1 , DataOut2 , DataOut3 , DataOut4 , DataOut5 , DataOut6 , DataOut7 , DataOut8 , DataOut9 , DataOut10 , DataOut11 , DataOut12 , DataOut13 , DataOut14 , DataOut15 , DataOut16 , DataOut17 , DataOut18 , DataOut19 , DataOut20 , DataOut21 , DataOut22 , DataOut23 , DataOut24 , DataOut25 , DataOut26 , DataOut27 , DataOut28 , DataOut29 , DataOut30 , DataOut31 , DataOut32 , DataOut33 , DataOut34 , DataOut35 , DataOut36 , DataOut37 , DataOut38 , DataOut39 , DataOut40 , DataOut41 , DataOut42 , DataOut43 , DataOut44 , DataOut45 , DataOut46 , DataOut47 , DataOut48 , DataOut49 , DataOut50 , DataOut51 , DataOut52 , DataOut53 , DataOut54 , DataOut55 , DataOut56 , DataOut57 , DataOut58 , DataOut59 , DataOut60 , DataOut61 , DataOut62 , DataOut63 , DataOut64 , DataOut65 , DataOut66 , DataOut67 , DataOut68 , DataOut69 , DataOut70 , DataOut71 , DataOut72 , DataOut73 , DataOut74 , DataOut75 , DataOut76 , DataOut77 , DataOut78 , DataOut79 , DataOut80 , DataOut81 , DataOut82 , DataOut83 , DataOut84 , DataOut85 , DataOut86 , DataOut87 , DataOut88 , DataOut89 , DataOut90 , DataOut91 , DataOut92 , DataOut93 , DataOut94 , DataOut95 , DataOut96 , DataOut97 , DataOut98 , DataOut99 , DataOut100 , DataOut101 , DataOut102 , DataOut103 , DataOut104 , DataOut105 , DataOut106 , DataOut107 , DataOut108 , DataOut109 , DataOut110 , DataOut111 , DataOut112 , DataOut113 , DataOut114 , DataOut115 , DataOut116 , DataOut117 , DataOut118 , DataOut119 , DataOut120 , DataOut121 , DataOut122 , DataOut123 , DataOut124 , DataOut125 , DataOut126 , DataOut127 , DataOut128 , DataOut129 , DataOut130 , DataOut131 , DataOut132 , DataOut133 , DataOut134 , DataOut135 , DataOut136 , DataOut137 , DataOut138 , DataOut139 , DataOut140 , DataOut141 , DataOut142 , DataOut143 , DataOut144 , DataOut145 , DataOut146 , DataOut147 , DataOut148 , DataOut149 , DataOut150 , DataOut151 , DataOut152 , DataOut153 , DataOut154 , DataOut155 , DataOut156 , DataOut157 , DataOut158 , DataOut159 , DataOut160 , DataOut161 , DataOut162 , DataOut163 , DataOut164 , DataOut165 , DataOut166 , DataOut167 , DataOut168 , DataOut169 , DataOut170 , DataOut171 , DataOut172 , DataOut173 , DataOut174 , DataOut175 , DataOut176 , DataOut177 , DataOut178 , DataOut179 , DataOut180 , DataOut181 , DataOut182 , DataOut183 , DataOut184 , DataOut185 , DataOut186 , DataOut187 , DataOut188 , DataOut189 , DataOut190 , DataOut191 , DataOut192 , DataOut193 , DataOut194 , DataOut195 , DataOut196 , DataOut197 , DataOut198 , DataOut199 , DataOut200 , DataOut201 , DataOut202 , DataOut203 , DataOut204 , DataOut205 , DataOut206 , DataOut207 , DataOut208 , DataOut209 , DataOut210 , DataOut211 , DataOut212 , DataOut213 , DataOut214 , DataOut215 , DataOut216 , DataOut217 , DataOut218 , DataOut219 , DataOut220 , DataOut221 , DataOut222 , DataOut223 , DataOut224 , DataOut225 , DataOut226 , DataOut227 , DataOut228 , DataOut229 , DataOut230 , DataOut231 , DataOut232 , DataOut233 , DataOut234 , DataOut235 , DataOut236 , DataOut237 , DataOut238 , DataOut239 , DataOut240 , DataOut241 , DataOut242 , DataOut243 , DataOut244 , DataOut245 , DataOut246 , DataOut247 , DataOut248 , DataOut249 , DataOut250 , DataOut251 , DataOut252 , DataOut253 , DataOut254 , DataOut255 , DataOut256 , DataOut257 , DataOut258 , DataOut259 , DataOut260 , DataOut261 , DataOut262 , DataOut263 , DataOut264 , DataOut265 , DataOut266 , DataOut267 , DataOut268 , DataOut269 , DataOut270 , DataOut271 , DataOut272 , DataOut273 , DataOut274 , DataOut275 , DataOut276 , DataOut277 , DataOut278 , DataOut279 , DataOut280 , DataOut281 , DataOut282 , DataOut283 , DataOut284 , DataOut285 , DataOut286 , DataOut287 , DataOut288 , DataOut289 , DataOut290 , DataOut291 , DataOut292 , DataOut293 , DataOut294 , DataOut295 , DataOut296 , DataOut297 , DataOut298 , DataOut299 , DataOut300 , DataOut301 , DataOut302 , DataOut303 , DataOut304 , DataOut305 , DataOut306 , DataOut307 , DataOut308 , DataOut309 , DataOut310 , DataOut311 , DataOut312 , DataOut313 , DataOut314 , DataOut315 , DataOut316 , DataOut317 , DataOut318 , DataOut319 , DataOut320 , DataOut321 , DataOut322 , DataOut323 , DataOut324 , DataOut325 , DataOut326 , DataOut327 , DataOut328 , DataOut329 , DataOut330 , DataOut331 , DataOut332 , DataOut333 , DataOut334 , DataOut335 , DataOut336 , DataOut337 , DataOut338 , DataOut339 , DataOut340 , DataOut341 , DataOut342 , DataOut343 , DataOut344 , DataOut345 , DataOut346 , DataOut347 , DataOut348 , DataOut349 , DataOut350 , DataOut351 , DataOut352 , DataOut353 , DataOut354 , DataOut355 , DataOut356 , DataOut357 , DataOut358 , DataOut359 , DataOut360 , DataOut361 , DataOut362 , DataOut363 , DataOut364 , DataOut365 , DataOut366 , DataOut367 , DataOut368 , DataOut369 , DataOut370 , DataOut371 , DataOut372 , DataOut373 , DataOut374 , DataOut375 , DataOut376 , DataOut377 , DataOut378 , DataOut379 , DataOut380 , DataOut381 , DataOut382 , DataOut383 , DataOut384 , DataOut385 , DataOut386 , DataOut387 , DataOut388 , DataOut389 , DataOut390 , DataOut391 , DataOut392 , DataOut393 , DataOut394 , DataOut395 , DataOut396 , DataOut397 , DataOut398 , DataOut399 , DataOut400 , DataOut401 , DataOut402 , DataOut403 , DataOut404 , DataOut405 , DataOut406 , DataOut407 , DataOut408 , DataOut409 , DataOut410 , DataOut411 , DataOut412 , DataOut413 , DataOut414 , DataOut415 , DataOut416 , DataOut417 , DataOut418 , DataOut419 , DataOut420 , DataOut421 , DataOut422 , DataOut423 , DataOut424 , DataOut425 , DataOut426 , DataOut427 , DataOut428 , DataOut429 , DataOut430 , DataOut431 , DataOut432 , DataOut433 , DataOut434 , DataOut435 , DataOut436 , DataOut437 , DataOut438 , DataOut439 , DataOut440 , DataOut441 , DataOut442 , DataOut443 , DataOut444 , DataOut445 , DataOut446 , DataOut447 , DataOut448 , DataOut449 , DataOut450 , DataOut451 , DataOut452 , DataOut453 , DataOut454 , DataOut455 , DataOut456 , DataOut457 , DataOut458 , DataOut459 , DataOut460 , DataOut461 , DataOut462 , DataOut463 , DataOut464 , DataOut465 , DataOut466 , DataOut467 , DataOut468 , DataOut469 , DataOut470 , DataOut471 , DataOut472 , DataOut473 , DataOut474 , DataOut475 , DataOut476 , DataOut477 , DataOut478 , DataOut479 , DataOut480 , DataOut481 , DataOut482 , DataOut483 , DataOut484 , DataOut485 , DataOut486 , DataOut487 , DataOut488 , DataOut489 , DataOut490 , DataOut491 , DataOut492 , DataOut493 , DataOut494 , DataOut495 , DataOut496 , DataOut497 , DataOut498 , DataOut499 , DataOut500 , DataOut501 , DataOut502 , DataOut503 , DataOut504 , DataOut505 , DataOut506 , DataOut507 , DataOut508 , DataOut509 , DataOut510 , DataOut511 , DataOut512 , DataOut513 , DataOut514 , DataOut515 , DataOut516 , DataOut517 , DataOut518 , DataOut519 , DataOut520 , DataOut521 , DataOut522 , DataOut523 , DataOut524 , DataOut525 , DataOut526 , DataOut527 , DataOut528 , DataOut529 , DataOut530 , DataOut531 , DataOut532 , DataOut533 , DataOut534 , DataOut535 , DataOut536 , DataOut537 , DataOut538 , DataOut539 , DataOut540 , DataOut541 , DataOut542 , DataOut543 , DataOut544 , DataOut545 , DataOut546 , DataOut547 , DataOut548 , DataOut549 , DataOut550 , DataOut551 , DataOut552 , DataOut553 , DataOut554 , DataOut555 , DataOut556 , DataOut557 , DataOut558 , DataOut559 , DataOut560 , DataOut561 , DataOut562 , DataOut563 , DataOut564 , DataOut565 , DataOut566 , DataOut567 , DataOut568 , DataOut569 , DataOut570 , DataOut571 , DataOut572 , DataOut573 , DataOut574 , DataOut575 , DataOut576 , DataOut577 , DataOut578 , DataOut579 , DataOut580 , DataOut581 , DataOut582 , DataOut583 , DataOut584 , DataOut585 , DataOut586 , DataOut587 , DataOut588 , DataOut589 , DataOut590 , DataOut591 , DataOut592 , DataOut593 , DataOut594 , DataOut595 , DataOut596 , DataOut597 , DataOut598 , DataOut599 , DataOut600 , DataOut601 , DataOut602 , DataOut603 , DataOut604 , DataOut605 , DataOut606 , DataOut607 , DataOut608 , DataOut609 , DataOut610 , DataOut611 , DataOut612 , DataOut613 , DataOut614 , DataOut615 , DataOut616 , DataOut617 , DataOut618 , DataOut619 , DataOut620 , DataOut621 , DataOut622 , DataOut623 , DataOut624 , DataOut625 , DataOut626 , DataOut627 , DataOut628 , DataOut629 , DataOut630 , DataOut631 , DataOut632 , DataOut633 , DataOut634 , DataOut635 , DataOut636 , DataOut637 , DataOut638 , DataOut639 , DataOut640 , DataOut641 , DataOut642 , DataOut643 , DataOut644 , DataOut645 , DataOut646 , DataOut647 , DataOut648 , DataOut649 , DataOut650 , DataOut651 , DataOut652 , DataOut653 , DataOut654 , DataOut655 , DataOut656 , DataOut657 , DataOut658 , DataOut659 , DataOut660 , DataOut661 , DataOut662 , DataOut663 , DataOut664 , DataOut665 , DataOut666 , DataOut667 , DataOut668 , DataOut669 , DataOut670 , DataOut671 , DataOut672 , DataOut673 , DataOut674 , DataOut675 , DataOut676 , DataOut677 , DataOut678 , DataOut679 , DataOut680 , DataOut681 , DataOut682 , DataOut683 , DataOut684 , DataOut685 , DataOut686 , DataOut687 , DataOut688 , DataOut689 , DataOut690 , DataOut691 , DataOut692 , DataOut693 , DataOut694 , DataOut695 , DataOut696 , DataOut697 , DataOut698 , DataOut699 , DataOut700 , DataOut701 , DataOut702 , DataOut703 , DataOut704 , DataOut705 , DataOut706 , DataOut707 , DataOut708 , DataOut709 , DataOut710 , DataOut711 , DataOut712 , DataOut713 , DataOut714 , DataOut715 , DataOut716 , DataOut717 , DataOut718 , DataOut719 , DataOut720 , DataOut721 , DataOut722 , DataOut723 , DataOut724 , DataOut725 , DataOut726 , DataOut727 , DataOut728 , DataOut729 , DataOut730 , DataOut731 , DataOut732 , DataOut733 , DataOut734 , DataOut735 , DataOut736 , DataOut737 , DataOut738 , DataOut739 , DataOut740 , DataOut741 , DataOut742 , DataOut743 , DataOut744 , DataOut745 , DataOut746 , DataOut747 , DataOut748 , DataOut749 , DataOut750 , DataOut751 , DataOut752 , DataOut753 , DataOut754 , DataOut755 , DataOut756 , DataOut757 , DataOut758 , DataOut759 , DataOut760 , DataOut761 , DataOut762 , DataOut763 , DataOut764 , DataOut765 , DataOut766 , DataOut767 , DataOut768 , DataOut769 , DataOut770 , DataOut771 , DataOut772 , DataOut773 , DataOut774 , DataOut775 , DataOut776 , DataOut777 , DataOut778 , DataOut779 , DataOut780 , DataOut781 , DataOut782 , DataOut783 ;
reg [65:0] DataOut784 = 66'b010011111111110000000000000000000000000000000000000000000000000000;
input Conv1LayerStart;
//output Conv1LayerFinish;


output MAX1LayerFinish;

output wire [65:0]  REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143; 
output wire [65:0]  REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143; 
output wire [65:0]  REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143; 
output wire [65:0]  REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143; 
 




//wire write2;
reg write2_1, write2_2, write2_3, write2_4, write2_5, write2_6, write2_7, write2_8, write2_9, write2_10, write2_11, write2_12, write2_13, write2_14, write2_15, write2_16, write2_17, write2_18, write2_19, write2_20, write2_21, write2_22, write2_23, write2_24, write2_25, write2_26, write2_27, write2_28, write2_29, write2_30, write2_31, write2_32, write2_33, write2_34, write2_35, write2_36, write2_37, write2_38, write2_39, write2_40, write2_41, write2_42, write2_43, write2_44, write2_45, write2_46, write2_47, write2_48, write2_49, write2_50, write2_51, write2_52, write2_53, write2_54, write2_55, write2_56, write2_57, write2_58, write2_59, write2_60, write2_61, write2_62, write2_63, write2_64, write2_65, write2_66, write2_67, write2_68, write2_69, write2_70, write2_71, write2_72, write2_73, write2_74, write2_75, write2_76, write2_77, write2_78, write2_79, write2_80, write2_81, write2_82, write2_83, write2_84, write2_85, write2_86, write2_87, write2_88, write2_89, write2_90, write2_91, write2_92, write2_93, write2_94, write2_95, write2_96, write2_97, write2_98, write2_99, write2_100, write2_101, write2_102, write2_103, write2_104, write2_105, write2_106, write2_107, write2_108, write2_109, write2_110, write2_111, write2_112, write2_113, write2_114, write2_115, write2_116, write2_117, write2_118, write2_119, write2_120, write2_121, write2_122, write2_123, write2_124, write2_125, write2_126, write2_127, write2_128, write2_129, write2_130, write2_131, write2_132, write2_133, write2_134, write2_135, write2_136, write2_137, write2_138, write2_139, write2_140, write2_141, write2_142, write2_143, write2_144;

wire  MAC_start, MAC_end;
wire [8:0] counter; 
wire [65:0]  ROMout1 , ROMout2 , ROMout3 , ROMout4;
wire [4:0]  address; 
wire [15:0] bigaddress;
wire [7:0] bigaddress340;


wire [65:0] Super_1_1_1_1 , Super_1_2_1_1 , Super_1_3_1_1 , Super_1_4_1_1 , Super_1_5_1_1 , Super_2_1_1_1 , Super_2_2_1_1 , Super_2_3_1_1 , Super_2_4_1_1 , Super_2_5_1_1 , Super_3_1_1_1 , Super_3_2_1_1 , Super_3_3_1_1 , Super_3_4_1_1 , Super_3_5_1_1 , Super_4_1_1_1 , Super_4_2_1_1 , Super_4_3_1_1 , Super_4_4_1_1 , Super_4_5_1_1 , Super_5_1_1_1 , Super_5_2_1_1 , Super_5_3_1_1 , Super_5_4_1_1 , Super_5_5_1_1 ;
wire [65:0] Super_1_1_1_2 , Super_1_2_1_2 , Super_1_3_1_2 , Super_1_4_1_2 , Super_1_5_1_2 , Super_2_1_1_2 , Super_2_2_1_2 , Super_2_3_1_2 , Super_2_4_1_2 , Super_2_5_1_2 , Super_3_1_1_2 , Super_3_2_1_2 , Super_3_3_1_2 , Super_3_4_1_2 , Super_3_5_1_2 , Super_4_1_1_2 , Super_4_2_1_2 , Super_4_3_1_2 , Super_4_4_1_2 , Super_4_5_1_2 , Super_5_1_1_2 , Super_5_2_1_2 , Super_5_3_1_2 , Super_5_4_1_2 , Super_5_5_1_2 ;
wire [65:0] Super_1_1_2_1 , Super_1_2_2_1 , Super_1_3_2_1 , Super_1_4_2_1 , Super_1_5_2_1 , Super_2_1_2_1 , Super_2_2_2_1 , Super_2_3_2_1 , Super_2_4_2_1 , Super_2_5_2_1 , Super_3_1_2_1 , Super_3_2_2_1 , Super_3_3_2_1 , Super_3_4_2_1 , Super_3_5_2_1 , Super_4_1_2_1 , Super_4_2_2_1 , Super_4_3_2_1 , Super_4_4_2_1 , Super_4_5_2_1 , Super_5_1_2_1 , Super_5_2_2_1 , Super_5_3_2_1 , Super_5_4_2_1 , Super_5_5_2_1 ;
wire [65:0] Super_1_1_2_2 , Super_1_2_2_2 , Super_1_3_2_2 , Super_1_4_2_2 , Super_1_5_2_2 , Super_2_1_2_2 , Super_2_2_2_2 , Super_2_3_2_2 , Super_2_4_2_2 , Super_2_5_2_2 , Super_3_1_2_2 , Super_3_2_2_2 , Super_3_3_2_2 , Super_3_4_2_2 , Super_3_5_2_2 , Super_4_1_2_2 , Super_4_2_2_2 , Super_4_3_2_2 , Super_4_4_2_2 , Super_4_5_2_2 , Super_5_1_2_2 , Super_5_2_2_2 , Super_5_3_2_2 , Super_5_4_2_2 , Super_5_5_2_2 ;





wire [65:0] MUXout1_1 , MUXout1_2 ;
wire [65:0] MUXout2_1 , MUXout2_2 ;




wire [65:0] MACout_F1_1_1  , MACout_F1_1_2  ,  MACout_F1_2_1  , MACout_F1_2_2  ;
wire [65:0] MACout_F2_1_1  , MACout_F2_1_2  ,  MACout_F2_2_1  , MACout_F2_2_2  ;
wire [65:0] MACout_F3_1_1  , MACout_F3_1_2  ,  MACout_F3_2_1  , MACout_F3_2_2  ;
wire [65:0] MACout_F4_1_1  , MACout_F4_1_2  ,  MACout_F4_2_1  , MACout_F4_2_2  ;


wire [65:0] RELUout_F1_1_1  , RELUout_F1_1_2    , RELUout_F1_2_1  , RELUout_F1_2_2  ;
wire [65:0] RELUout_F2_1_1  , RELUout_F2_1_2    , RELUout_F2_2_1  , RELUout_F2_2_2  ;
wire [65:0] RELUout_F3_1_1  , RELUout_F3_1_2    , RELUout_F3_2_1  , RELUout_F3_2_2  ;
wire [65:0] RELUout_F4_1_1  , RELUout_F4_1_2    , RELUout_F4_2_1  , RELUout_F4_2_2  ;


/* 
output wire [65:0] Final_1_F1_1_1  , Final_1_F1_1_2  , Final_1_F1_2_1  , Final_1_F1_2_2  ;
output wire [65:0] Final_1_F2_1_1  , Final_1_F2_1_2  , Final_1_F2_2_1  , Final_1_F2_2_2  ;
output wire [65:0] Final_1_F3_1_1  , Final_1_F3_1_2  , Final_1_F3_2_1  , Final_1_F3_2_2  ;
output wire [65:0] Final_1_F4_1_1  , Final_1_F4_1_2  , Final_1_F4_2_1  , Final_1_F4_2_2  ;
output wire [65:0] Final_2_F1_1_1  , Final_2_F1_1_2  , Final_2_F1_2_1  , Final_2_F1_2_2  ;
output wire [65:0] Final_2_F2_1_1  , Final_2_F2_1_2  , Final_2_F2_2_1  , Final_2_F2_2_2  ;
output wire [65:0] Final_2_F3_1_1  , Final_2_F3_1_2  , Final_2_F3_2_1  , Final_2_F3_2_2  ;
output wire [65:0] Final_2_F4_1_1  , Final_2_F4_1_2  , Final_2_F4_2_1  , Final_2_F4_2_2  ;
output wire [65:0] Final_3_F1_1_1  , Final_3_F1_1_2  , Final_3_F1_2_1  , Final_3_F1_2_2  ;
output wire [65:0] Final_3_F2_1_1  , Final_3_F2_1_2  , Final_3_F2_2_1  , Final_3_F2_2_2  ;
output wire [65:0] Final_3_F3_1_1  , Final_3_F3_1_2  , Final_3_F3_2_1  , Final_3_F3_2_2  ;
output wire [65:0] Final_3_F4_1_1  , Final_3_F4_1_2  , Final_3_F4_2_1  , Final_3_F4_2_2  ;
output wire [65:0] Final_4_F1_1_1  , Final_4_F1_1_2  , Final_4_F1_2_1  , Final_4_F1_2_2  ;
output wire [65:0] Final_4_F2_1_1  , Final_4_F2_1_2  , Final_4_F2_2_1  , Final_4_F2_2_2  ;
output wire [65:0] Final_4_F3_1_1  , Final_4_F3_1_2  , Final_4_F3_2_1  , Final_4_F3_2_2  ;
output wire [65:0] Final_4_F4_1_1  , Final_4_F4_1_2  , Final_4_F4_2_1  , Final_4_F4_2_2  ;
output wire [65:0] Final_5_F1_1_1  , Final_5_F1_1_2  , Final_5_F1_2_1  , Final_5_F1_2_2  ;
output wire [65:0] Final_5_F2_1_1  , Final_5_F2_1_2  , Final_5_F2_2_1  , Final_5_F2_2_2  ;
output wire [65:0] Final_5_F3_1_1  , Final_5_F3_1_2  , Final_5_F3_2_1  , Final_5_F3_2_2  ;
output wire [65:0] Final_5_F4_1_1  , Final_5_F4_1_2  , Final_5_F4_2_1  , Final_5_F4_2_2  ;
output wire [65:0] Final_6_F1_1_1  , Final_6_F1_1_2  , Final_6_F1_2_1  , Final_6_F1_2_2  ;
output wire [65:0] Final_6_F2_1_1  , Final_6_F2_1_2  , Final_6_F2_2_1  , Final_6_F2_2_2  ;
output wire [65:0] Final_6_F3_1_1  , Final_6_F3_1_2  , Final_6_F3_2_1  , Final_6_F3_2_2  ;
output wire [65:0] Final_6_F4_1_1  , Final_6_F4_1_2  , Final_6_F4_2_1  , Final_6_F4_2_2  ;
output wire [65:0] Final_7_F1_1_1  , Final_7_F1_1_2  , Final_7_F1_2_1  , Final_7_F1_2_2  ;
output wire [65:0] Final_7_F2_1_1  , Final_7_F2_1_2  , Final_7_F2_2_1  , Final_7_F2_2_2  ;
output wire [65:0] Final_7_F3_1_1  , Final_7_F3_1_2  , Final_7_F3_2_1  , Final_7_F3_2_2  ;
output wire [65:0] Final_7_F4_1_1  , Final_7_F4_1_2  , Final_7_F4_2_1  , Final_7_F4_2_2  ;
output wire [65:0] Final_8_F1_1_1  , Final_8_F1_1_2  , Final_8_F1_2_1  , Final_8_F1_2_2  ;
output wire [65:0] Final_8_F2_1_1  , Final_8_F2_1_2  , Final_8_F2_2_1  , Final_8_F2_2_2  ;
output wire [65:0] Final_8_F3_1_1  , Final_8_F3_1_2  , Final_8_F3_2_1  , Final_8_F3_2_2  ;
output wire [65:0] Final_8_F4_1_1  , Final_8_F4_1_2  , Final_8_F4_2_1  , Final_8_F4_2_2  ;
output wire [65:0] Final_9_F1_1_1  , Final_9_F1_1_2  , Final_9_F1_2_1  , Final_9_F1_2_2  ;
output wire [65:0] Final_9_F2_1_1  , Final_9_F2_1_2  , Final_9_F2_2_1  , Final_9_F2_2_2  ;
output wire [65:0] Final_9_F3_1_1  , Final_9_F3_1_2  , Final_9_F3_2_1  , Final_9_F3_2_2  ;
output wire [65:0] Final_9_F4_1_1  , Final_9_F4_1_2  , Final_9_F4_2_1  , Final_9_F4_2_2  ;
output wire [65:0] Final_10_F1_1_1  , Final_10_F1_1_2  , Final_10_F1_2_1  , Final_10_F1_2_2  ;
output wire [65:0] Final_10_F2_1_1  , Final_10_F2_1_2  , Final_10_F2_2_1  , Final_10_F2_2_2  ;
output wire [65:0] Final_10_F3_1_1  , Final_10_F3_1_2  , Final_10_F3_2_1  , Final_10_F3_2_2  ;
output wire [65:0] Final_10_F4_1_1  , Final_10_F4_1_2  , Final_10_F4_2_1  , Final_10_F4_2_2  ;
output wire [65:0] Final_11_F1_1_1  , Final_11_F1_1_2  , Final_11_F1_2_1  , Final_11_F1_2_2  ;
output wire [65:0] Final_11_F2_1_1  , Final_11_F2_1_2  , Final_11_F2_2_1  , Final_11_F2_2_2  ;
output wire [65:0] Final_11_F3_1_1  , Final_11_F3_1_2  , Final_11_F3_2_1  , Final_11_F3_2_2  ;
output wire [65:0] Final_11_F4_1_1  , Final_11_F4_1_2  , Final_11_F4_2_1  , Final_11_F4_2_2  ;
output wire [65:0] Final_12_F1_1_1  , Final_12_F1_1_2  , Final_12_F1_2_1  , Final_12_F1_2_2  ;
output wire [65:0] Final_12_F2_1_1  , Final_12_F2_1_2  , Final_12_F2_2_1  , Final_12_F2_2_2  ;
output wire [65:0] Final_12_F3_1_1  , Final_12_F3_1_2  , Final_12_F3_2_1  , Final_12_F3_2_2  ;
output wire [65:0] Final_12_F4_1_1  , Final_12_F4_1_2  , Final_12_F4_2_1  , Final_12_F4_2_2  ;
output wire [65:0] Final_13_F1_1_1  , Final_13_F1_1_2  , Final_13_F1_2_1  , Final_13_F1_2_2  ;
output wire [65:0] Final_13_F2_1_1  , Final_13_F2_1_2  , Final_13_F2_2_1  , Final_13_F2_2_2  ;
output wire [65:0] Final_13_F3_1_1  , Final_13_F3_1_2  , Final_13_F3_2_1  , Final_13_F3_2_2  ;
output wire [65:0] Final_13_F4_1_1  , Final_13_F4_1_2  , Final_13_F4_2_1  , Final_13_F4_2_2  ;
output wire [65:0] Final_14_F1_1_1  , Final_14_F1_1_2  , Final_14_F1_2_1  , Final_14_F1_2_2  ;
output wire [65:0] Final_14_F2_1_1  , Final_14_F2_1_2  , Final_14_F2_2_1  , Final_14_F2_2_2  ;
output wire [65:0] Final_14_F3_1_1  , Final_14_F3_1_2  , Final_14_F3_2_1  , Final_14_F3_2_2  ;
output wire [65:0] Final_14_F4_1_1  , Final_14_F4_1_2  , Final_14_F4_2_1  , Final_14_F4_2_2  ;
output wire [65:0] Final_15_F1_1_1  , Final_15_F1_1_2  , Final_15_F1_2_1  , Final_15_F1_2_2  ;
output wire [65:0] Final_15_F2_1_1  , Final_15_F2_1_2  , Final_15_F2_2_1  , Final_15_F2_2_2  ;
output wire [65:0] Final_15_F3_1_1  , Final_15_F3_1_2  , Final_15_F3_2_1  , Final_15_F3_2_2  ;
output wire [65:0] Final_15_F4_1_1  , Final_15_F4_1_2  , Final_15_F4_2_1  , Final_15_F4_2_2  ;
output wire [65:0] Final_16_F1_1_1  , Final_16_F1_1_2  , Final_16_F1_2_1  , Final_16_F1_2_2  ;
output wire [65:0] Final_16_F2_1_1  , Final_16_F2_1_2  , Final_16_F2_2_1  , Final_16_F2_2_2  ;
output wire [65:0] Final_16_F3_1_1  , Final_16_F3_1_2  , Final_16_F3_2_1  , Final_16_F3_2_2  ;
output wire [65:0] Final_16_F4_1_1  , Final_16_F4_1_2  , Final_16_F4_2_1  , Final_16_F4_2_2  ;
output wire [65:0] Final_17_F1_1_1  , Final_17_F1_1_2  , Final_17_F1_2_1  , Final_17_F1_2_2  ;
output wire [65:0] Final_17_F2_1_1  , Final_17_F2_1_2  , Final_17_F2_2_1  , Final_17_F2_2_2  ;
output wire [65:0] Final_17_F3_1_1  , Final_17_F3_1_2  , Final_17_F3_2_1  , Final_17_F3_2_2  ;
output wire [65:0] Final_17_F4_1_1  , Final_17_F4_1_2  , Final_17_F4_2_1  , Final_17_F4_2_2  ;
output wire [65:0] Final_18_F1_1_1  , Final_18_F1_1_2  , Final_18_F1_2_1  , Final_18_F1_2_2  ;
output wire [65:0] Final_18_F2_1_1  , Final_18_F2_1_2  , Final_18_F2_2_1  , Final_18_F2_2_2  ;
output wire [65:0] Final_18_F3_1_1  , Final_18_F3_1_2  , Final_18_F3_2_1  , Final_18_F3_2_2  ;
output wire [65:0] Final_18_F4_1_1  , Final_18_F4_1_2  , Final_18_F4_2_1  , Final_18_F4_2_2  ;
output wire [65:0] Final_19_F1_1_1  , Final_19_F1_1_2  , Final_19_F1_2_1  , Final_19_F1_2_2  ;
output wire [65:0] Final_19_F2_1_1  , Final_19_F2_1_2  , Final_19_F2_2_1  , Final_19_F2_2_2  ;
output wire [65:0] Final_19_F3_1_1  , Final_19_F3_1_2  , Final_19_F3_2_1  , Final_19_F3_2_2  ;
output wire [65:0] Final_19_F4_1_1  , Final_19_F4_1_2  , Final_19_F4_2_1  , Final_19_F4_2_2  ;
output wire [65:0] Final_20_F1_1_1  , Final_20_F1_1_2  , Final_20_F1_2_1  , Final_20_F1_2_2  ;
output wire [65:0] Final_20_F2_1_1  , Final_20_F2_1_2  , Final_20_F2_2_1  , Final_20_F2_2_2  ;
output wire [65:0] Final_20_F3_1_1  , Final_20_F3_1_2  , Final_20_F3_2_1  , Final_20_F3_2_2  ;
output wire [65:0] Final_20_F4_1_1  , Final_20_F4_1_2  , Final_20_F4_2_1  , Final_20_F4_2_2  ;
output wire [65:0] Final_21_F1_1_1  , Final_21_F1_1_2  , Final_21_F1_2_1  , Final_21_F1_2_2  ;
output wire [65:0] Final_21_F2_1_1  , Final_21_F2_1_2  , Final_21_F2_2_1  , Final_21_F2_2_2  ;
output wire [65:0] Final_21_F3_1_1  , Final_21_F3_1_2  , Final_21_F3_2_1  , Final_21_F3_2_2  ;
output wire [65:0] Final_21_F4_1_1  , Final_21_F4_1_2  , Final_21_F4_2_1  , Final_21_F4_2_2  ;
output wire [65:0] Final_22_F1_1_1  , Final_22_F1_1_2  , Final_22_F1_2_1  , Final_22_F1_2_2  ;
output wire [65:0] Final_22_F2_1_1  , Final_22_F2_1_2  , Final_22_F2_2_1  , Final_22_F2_2_2  ;
output wire [65:0] Final_22_F3_1_1  , Final_22_F3_1_2  , Final_22_F3_2_1  , Final_22_F3_2_2  ;
output wire [65:0] Final_22_F4_1_1  , Final_22_F4_1_2  , Final_22_F4_2_1  , Final_22_F4_2_2  ;
output wire [65:0] Final_23_F1_1_1  , Final_23_F1_1_2  , Final_23_F1_2_1  , Final_23_F1_2_2  ;
output wire [65:0] Final_23_F2_1_1  , Final_23_F2_1_2  , Final_23_F2_2_1  , Final_23_F2_2_2  ;
output wire [65:0] Final_23_F3_1_1  , Final_23_F3_1_2  , Final_23_F3_2_1  , Final_23_F3_2_2  ;
output wire [65:0] Final_23_F4_1_1  , Final_23_F4_1_2  , Final_23_F4_2_1  , Final_23_F4_2_2  ;
output wire [65:0] Final_24_F1_1_1  , Final_24_F1_1_2  , Final_24_F1_2_1  , Final_24_F1_2_2  ;
output wire [65:0] Final_24_F2_1_1  , Final_24_F2_1_2  , Final_24_F2_2_1  , Final_24_F2_2_2  ;
output wire [65:0] Final_24_F3_1_1  , Final_24_F3_1_2  , Final_24_F3_2_1  , Final_24_F3_2_2  ;
output wire [65:0] Final_24_F4_1_1  , Final_24_F4_1_2  , Final_24_F4_2_1  , Final_24_F4_2_2  ;
output wire [65:0] Final_25_F1_1_1  , Final_25_F1_1_2  , Final_25_F1_2_1  , Final_25_F1_2_2  ;
output wire [65:0] Final_25_F2_1_1  , Final_25_F2_1_2  , Final_25_F2_2_1  , Final_25_F2_2_2  ;
output wire [65:0] Final_25_F3_1_1  , Final_25_F3_1_2  , Final_25_F3_2_1  , Final_25_F3_2_2  ;
output wire [65:0] Final_25_F4_1_1  , Final_25_F4_1_2  , Final_25_F4_2_1  , Final_25_F4_2_2  ;
output wire [65:0] Final_26_F1_1_1  , Final_26_F1_1_2  , Final_26_F1_2_1  , Final_26_F1_2_2  ;
output wire [65:0] Final_26_F2_1_1  , Final_26_F2_1_2  , Final_26_F2_2_1  , Final_26_F2_2_2  ;
output wire [65:0] Final_26_F3_1_1  , Final_26_F3_1_2  , Final_26_F3_2_1  , Final_26_F3_2_2  ;
output wire [65:0] Final_26_F4_1_1  , Final_26_F4_1_2  , Final_26_F4_2_1  , Final_26_F4_2_2  ;
output wire [65:0] Final_27_F1_1_1  , Final_27_F1_1_2  , Final_27_F1_2_1  , Final_27_F1_2_2  ;
output wire [65:0] Final_27_F2_1_1  , Final_27_F2_1_2  , Final_27_F2_2_1  , Final_27_F2_2_2  ;
output wire [65:0] Final_27_F3_1_1  , Final_27_F3_1_2  , Final_27_F3_2_1  , Final_27_F3_2_2  ;
output wire [65:0] Final_27_F4_1_1  , Final_27_F4_1_2  , Final_27_F4_2_1  , Final_27_F4_2_2  ;
output wire [65:0] Final_28_F1_1_1  , Final_28_F1_1_2  , Final_28_F1_2_1  , Final_28_F1_2_2  ;
output wire [65:0] Final_28_F2_1_1  , Final_28_F2_1_2  , Final_28_F2_2_1  , Final_28_F2_2_2  ;
output wire [65:0] Final_28_F3_1_1  , Final_28_F3_1_2  , Final_28_F3_2_1  , Final_28_F3_2_2  ;
output wire [65:0] Final_28_F4_1_1  , Final_28_F4_1_2  , Final_28_F4_2_1  , Final_28_F4_2_2  ;
output wire [65:0] Final_29_F1_1_1  , Final_29_F1_1_2  , Final_29_F1_2_1  , Final_29_F1_2_2  ;
output wire [65:0] Final_29_F2_1_1  , Final_29_F2_1_2  , Final_29_F2_2_1  , Final_29_F2_2_2  ;
output wire [65:0] Final_29_F3_1_1  , Final_29_F3_1_2  , Final_29_F3_2_1  , Final_29_F3_2_2  ;
output wire [65:0] Final_29_F4_1_1  , Final_29_F4_1_2  , Final_29_F4_2_1  , Final_29_F4_2_2  ;
output wire [65:0] Final_30_F1_1_1  , Final_30_F1_1_2  , Final_30_F1_2_1  , Final_30_F1_2_2  ;
output wire [65:0] Final_30_F2_1_1  , Final_30_F2_1_2  , Final_30_F2_2_1  , Final_30_F2_2_2  ;
output wire [65:0] Final_30_F3_1_1  , Final_30_F3_1_2  , Final_30_F3_2_1  , Final_30_F3_2_2  ;
output wire [65:0] Final_30_F4_1_1  , Final_30_F4_1_2  , Final_30_F4_2_1  , Final_30_F4_2_2  ;
output wire [65:0] Final_31_F1_1_1  , Final_31_F1_1_2  , Final_31_F1_2_1  , Final_31_F1_2_2  ;
output wire [65:0] Final_31_F2_1_1  , Final_31_F2_1_2  , Final_31_F2_2_1  , Final_31_F2_2_2  ;
output wire [65:0] Final_31_F3_1_1  , Final_31_F3_1_2  , Final_31_F3_2_1  , Final_31_F3_2_2  ;
output wire [65:0] Final_31_F4_1_1  , Final_31_F4_1_2  , Final_31_F4_2_1  , Final_31_F4_2_2  ;
output wire [65:0] Final_32_F1_1_1  , Final_32_F1_1_2  , Final_32_F1_2_1  , Final_32_F1_2_2  ;
output wire [65:0] Final_32_F2_1_1  , Final_32_F2_1_2  , Final_32_F2_2_1  , Final_32_F2_2_2  ;
output wire [65:0] Final_32_F3_1_1  , Final_32_F3_1_2  , Final_32_F3_2_1  , Final_32_F3_2_2  ;
output wire [65:0] Final_32_F4_1_1  , Final_32_F4_1_2  , Final_32_F4_2_1  , Final_32_F4_2_2  ;
output wire [65:0] Final_33_F1_1_1  , Final_33_F1_1_2  , Final_33_F1_2_1  , Final_33_F1_2_2  ;
output wire [65:0] Final_33_F2_1_1  , Final_33_F2_1_2  , Final_33_F2_2_1  , Final_33_F2_2_2  ;
output wire [65:0] Final_33_F3_1_1  , Final_33_F3_1_2  , Final_33_F3_2_1  , Final_33_F3_2_2  ;
output wire [65:0] Final_33_F4_1_1  , Final_33_F4_1_2  , Final_33_F4_2_1  , Final_33_F4_2_2  ;
output wire [65:0] Final_34_F1_1_1  , Final_34_F1_1_2  , Final_34_F1_2_1  , Final_34_F1_2_2  ;
output wire [65:0] Final_34_F2_1_1  , Final_34_F2_1_2  , Final_34_F2_2_1  , Final_34_F2_2_2  ;
output wire [65:0] Final_34_F3_1_1  , Final_34_F3_1_2  , Final_34_F3_2_1  , Final_34_F3_2_2  ;
output wire [65:0] Final_34_F4_1_1  , Final_34_F4_1_2  , Final_34_F4_2_1  , Final_34_F4_2_2  ;
output wire [65:0] Final_35_F1_1_1  , Final_35_F1_1_2  , Final_35_F1_2_1  , Final_35_F1_2_2  ;
output wire [65:0] Final_35_F2_1_1  , Final_35_F2_1_2  , Final_35_F2_2_1  , Final_35_F2_2_2  ;
output wire [65:0] Final_35_F3_1_1  , Final_35_F3_1_2  , Final_35_F3_2_1  , Final_35_F3_2_2  ;
output wire [65:0] Final_35_F4_1_1  , Final_35_F4_1_2  , Final_35_F4_2_1  , Final_35_F4_2_2  ;
output wire [65:0] Final_36_F1_1_1  , Final_36_F1_1_2  , Final_36_F1_2_1  , Final_36_F1_2_2  ;
output wire [65:0] Final_36_F2_1_1  , Final_36_F2_1_2  , Final_36_F2_2_1  , Final_36_F2_2_2  ;
output wire [65:0] Final_36_F3_1_1  , Final_36_F3_1_2  , Final_36_F3_2_1  , Final_36_F3_2_2  ;
output wire [65:0] Final_36_F4_1_1  , Final_36_F4_1_2  , Final_36_F4_2_1  , Final_36_F4_2_2  ;
output wire [65:0] Final_37_F1_1_1  , Final_37_F1_1_2  , Final_37_F1_2_1  , Final_37_F1_2_2  ;
output wire [65:0] Final_37_F2_1_1  , Final_37_F2_1_2  , Final_37_F2_2_1  , Final_37_F2_2_2  ;
output wire [65:0] Final_37_F3_1_1  , Final_37_F3_1_2  , Final_37_F3_2_1  , Final_37_F3_2_2  ;
output wire [65:0] Final_37_F4_1_1  , Final_37_F4_1_2  , Final_37_F4_2_1  , Final_37_F4_2_2  ;
output wire [65:0] Final_38_F1_1_1  , Final_38_F1_1_2  , Final_38_F1_2_1  , Final_38_F1_2_2  ;
output wire [65:0] Final_38_F2_1_1  , Final_38_F2_1_2  , Final_38_F2_2_1  , Final_38_F2_2_2  ;
output wire [65:0] Final_38_F3_1_1  , Final_38_F3_1_2  , Final_38_F3_2_1  , Final_38_F3_2_2  ;
output wire [65:0] Final_38_F4_1_1  , Final_38_F4_1_2  , Final_38_F4_2_1  , Final_38_F4_2_2  ;
output wire [65:0] Final_39_F1_1_1  , Final_39_F1_1_2  , Final_39_F1_2_1  , Final_39_F1_2_2  ;
output wire [65:0] Final_39_F2_1_1  , Final_39_F2_1_2  , Final_39_F2_2_1  , Final_39_F2_2_2  ;
output wire [65:0] Final_39_F3_1_1  , Final_39_F3_1_2  , Final_39_F3_2_1  , Final_39_F3_2_2  ;
output wire [65:0] Final_39_F4_1_1  , Final_39_F4_1_2  , Final_39_F4_2_1  , Final_39_F4_2_2  ;
output wire [65:0] Final_40_F1_1_1  , Final_40_F1_1_2  , Final_40_F1_2_1  , Final_40_F1_2_2  ;
output wire [65:0] Final_40_F2_1_1  , Final_40_F2_1_2  , Final_40_F2_2_1  , Final_40_F2_2_2  ;
output wire [65:0] Final_40_F3_1_1  , Final_40_F3_1_2  , Final_40_F3_2_1  , Final_40_F3_2_2  ;
output wire [65:0] Final_40_F4_1_1  , Final_40_F4_1_2  , Final_40_F4_2_1  , Final_40_F4_2_2  ;
output wire [65:0] Final_41_F1_1_1  , Final_41_F1_1_2  , Final_41_F1_2_1  , Final_41_F1_2_2  ;
output wire [65:0] Final_41_F2_1_1  , Final_41_F2_1_2  , Final_41_F2_2_1  , Final_41_F2_2_2  ;
output wire [65:0] Final_41_F3_1_1  , Final_41_F3_1_2  , Final_41_F3_2_1  , Final_41_F3_2_2  ;
output wire [65:0] Final_41_F4_1_1  , Final_41_F4_1_2  , Final_41_F4_2_1  , Final_41_F4_2_2  ;
output wire [65:0] Final_42_F1_1_1  , Final_42_F1_1_2  , Final_42_F1_2_1  , Final_42_F1_2_2  ;
output wire [65:0] Final_42_F2_1_1  , Final_42_F2_1_2  , Final_42_F2_2_1  , Final_42_F2_2_2  ;
output wire [65:0] Final_42_F3_1_1  , Final_42_F3_1_2  , Final_42_F3_2_1  , Final_42_F3_2_2  ;
output wire [65:0] Final_42_F4_1_1  , Final_42_F4_1_2  , Final_42_F4_2_1  , Final_42_F4_2_2  ;
output wire [65:0] Final_43_F1_1_1  , Final_43_F1_1_2  , Final_43_F1_2_1  , Final_43_F1_2_2  ;
output wire [65:0] Final_43_F2_1_1  , Final_43_F2_1_2  , Final_43_F2_2_1  , Final_43_F2_2_2  ;
output wire [65:0] Final_43_F3_1_1  , Final_43_F3_1_2  , Final_43_F3_2_1  , Final_43_F3_2_2  ;
output wire [65:0] Final_43_F4_1_1  , Final_43_F4_1_2  , Final_43_F4_2_1  , Final_43_F4_2_2  ;
output wire [65:0] Final_44_F1_1_1  , Final_44_F1_1_2  , Final_44_F1_2_1  , Final_44_F1_2_2  ;
output wire [65:0] Final_44_F2_1_1  , Final_44_F2_1_2  , Final_44_F2_2_1  , Final_44_F2_2_2  ;
output wire [65:0] Final_44_F3_1_1  , Final_44_F3_1_2  , Final_44_F3_2_1  , Final_44_F3_2_2  ;
output wire [65:0] Final_44_F4_1_1  , Final_44_F4_1_2  , Final_44_F4_2_1  , Final_44_F4_2_2  ;
output wire [65:0] Final_45_F1_1_1  , Final_45_F1_1_2  , Final_45_F1_2_1  , Final_45_F1_2_2  ;
output wire [65:0] Final_45_F2_1_1  , Final_45_F2_1_2  , Final_45_F2_2_1  , Final_45_F2_2_2  ;
output wire [65:0] Final_45_F3_1_1  , Final_45_F3_1_2  , Final_45_F3_2_1  , Final_45_F3_2_2  ;
output wire [65:0] Final_45_F4_1_1  , Final_45_F4_1_2  , Final_45_F4_2_1  , Final_45_F4_2_2  ;
output wire [65:0] Final_46_F1_1_1  , Final_46_F1_1_2  , Final_46_F1_2_1  , Final_46_F1_2_2  ;
output wire [65:0] Final_46_F2_1_1  , Final_46_F2_1_2  , Final_46_F2_2_1  , Final_46_F2_2_2  ;
output wire [65:0] Final_46_F3_1_1  , Final_46_F3_1_2  , Final_46_F3_2_1  , Final_46_F3_2_2  ;
output wire [65:0] Final_46_F4_1_1  , Final_46_F4_1_2  , Final_46_F4_2_1  , Final_46_F4_2_2  ;
output wire [65:0] Final_47_F1_1_1  , Final_47_F1_1_2  , Final_47_F1_2_1  , Final_47_F1_2_2  ;
output wire [65:0] Final_47_F2_1_1  , Final_47_F2_1_2  , Final_47_F2_2_1  , Final_47_F2_2_2  ;
output wire [65:0] Final_47_F3_1_1  , Final_47_F3_1_2  , Final_47_F3_2_1  , Final_47_F3_2_2  ;
output wire [65:0] Final_47_F4_1_1  , Final_47_F4_1_2  , Final_47_F4_2_1  , Final_47_F4_2_2  ;
output wire [65:0] Final_48_F1_1_1  , Final_48_F1_1_2  , Final_48_F1_2_1  , Final_48_F1_2_2  ;
output wire [65:0] Final_48_F2_1_1  , Final_48_F2_1_2  , Final_48_F2_2_1  , Final_48_F2_2_2  ;
output wire [65:0] Final_48_F3_1_1  , Final_48_F3_1_2  , Final_48_F3_2_1  , Final_48_F3_2_2  ;
output wire [65:0] Final_48_F4_1_1  , Final_48_F4_1_2  , Final_48_F4_2_1  , Final_48_F4_2_2  ;
output wire [65:0] Final_49_F1_1_1  , Final_49_F1_1_2  , Final_49_F1_2_1  , Final_49_F1_2_2  ;
output wire [65:0] Final_49_F2_1_1  , Final_49_F2_1_2  , Final_49_F2_2_1  , Final_49_F2_2_2  ;
output wire [65:0] Final_49_F3_1_1  , Final_49_F3_1_2  , Final_49_F3_2_1  , Final_49_F3_2_2  ;
output wire [65:0] Final_49_F4_1_1  , Final_49_F4_1_2  , Final_49_F4_2_1  , Final_49_F4_2_2  ;
output wire [65:0] Final_50_F1_1_1  , Final_50_F1_1_2  , Final_50_F1_2_1  , Final_50_F1_2_2  ;
output wire [65:0] Final_50_F2_1_1  , Final_50_F2_1_2  , Final_50_F2_2_1  , Final_50_F2_2_2  ;
output wire [65:0] Final_50_F3_1_1  , Final_50_F3_1_2  , Final_50_F3_2_1  , Final_50_F3_2_2  ;
output wire [65:0] Final_50_F4_1_1  , Final_50_F4_1_2  , Final_50_F4_2_1  , Final_50_F4_2_2  ;
output wire [65:0] Final_51_F1_1_1  , Final_51_F1_1_2  , Final_51_F1_2_1  , Final_51_F1_2_2  ;
output wire [65:0] Final_51_F2_1_1  , Final_51_F2_1_2  , Final_51_F2_2_1  , Final_51_F2_2_2  ;
output wire [65:0] Final_51_F3_1_1  , Final_51_F3_1_2  , Final_51_F3_2_1  , Final_51_F3_2_2  ;
output wire [65:0] Final_51_F4_1_1  , Final_51_F4_1_2  , Final_51_F4_2_1  , Final_51_F4_2_2  ;
output wire [65:0] Final_52_F1_1_1  , Final_52_F1_1_2  , Final_52_F1_2_1  , Final_52_F1_2_2  ;
output wire [65:0] Final_52_F2_1_1  , Final_52_F2_1_2  , Final_52_F2_2_1  , Final_52_F2_2_2  ;
output wire [65:0] Final_52_F3_1_1  , Final_52_F3_1_2  , Final_52_F3_2_1  , Final_52_F3_2_2  ;
output wire [65:0] Final_52_F4_1_1  , Final_52_F4_1_2  , Final_52_F4_2_1  , Final_52_F4_2_2  ;
output wire [65:0] Final_53_F1_1_1  , Final_53_F1_1_2  , Final_53_F1_2_1  , Final_53_F1_2_2  ;
output wire [65:0] Final_53_F2_1_1  , Final_53_F2_1_2  , Final_53_F2_2_1  , Final_53_F2_2_2  ;
output wire [65:0] Final_53_F3_1_1  , Final_53_F3_1_2  , Final_53_F3_2_1  , Final_53_F3_2_2  ;
output wire [65:0] Final_53_F4_1_1  , Final_53_F4_1_2  , Final_53_F4_2_1  , Final_53_F4_2_2  ;
output wire [65:0] Final_54_F1_1_1  , Final_54_F1_1_2  , Final_54_F1_2_1  , Final_54_F1_2_2  ;
output wire [65:0] Final_54_F2_1_1  , Final_54_F2_1_2  , Final_54_F2_2_1  , Final_54_F2_2_2  ;
output wire [65:0] Final_54_F3_1_1  , Final_54_F3_1_2  , Final_54_F3_2_1  , Final_54_F3_2_2  ;
output wire [65:0] Final_54_F4_1_1  , Final_54_F4_1_2  , Final_54_F4_2_1  , Final_54_F4_2_2  ;
output wire [65:0] Final_55_F1_1_1  , Final_55_F1_1_2  , Final_55_F1_2_1  , Final_55_F1_2_2  ;
output wire [65:0] Final_55_F2_1_1  , Final_55_F2_1_2  , Final_55_F2_2_1  , Final_55_F2_2_2  ;
output wire [65:0] Final_55_F3_1_1  , Final_55_F3_1_2  , Final_55_F3_2_1  , Final_55_F3_2_2  ;
output wire [65:0] Final_55_F4_1_1  , Final_55_F4_1_2  , Final_55_F4_2_1  , Final_55_F4_2_2  ;
output wire [65:0] Final_56_F1_1_1  , Final_56_F1_1_2  , Final_56_F1_2_1  , Final_56_F1_2_2  ;
output wire [65:0] Final_56_F2_1_1  , Final_56_F2_1_2  , Final_56_F2_2_1  , Final_56_F2_2_2  ;
output wire [65:0] Final_56_F3_1_1  , Final_56_F3_1_2  , Final_56_F3_2_1  , Final_56_F3_2_2  ;
output wire [65:0] Final_56_F4_1_1  , Final_56_F4_1_2  , Final_56_F4_2_1  , Final_56_F4_2_2  ;
output wire [65:0] Final_57_F1_1_1  , Final_57_F1_1_2  , Final_57_F1_2_1  , Final_57_F1_2_2  ;
output wire [65:0] Final_57_F2_1_1  , Final_57_F2_1_2  , Final_57_F2_2_1  , Final_57_F2_2_2  ;
output wire [65:0] Final_57_F3_1_1  , Final_57_F3_1_2  , Final_57_F3_2_1  , Final_57_F3_2_2  ;
output wire [65:0] Final_57_F4_1_1  , Final_57_F4_1_2  , Final_57_F4_2_1  , Final_57_F4_2_2  ;
output wire [65:0] Final_58_F1_1_1  , Final_58_F1_1_2  , Final_58_F1_2_1  , Final_58_F1_2_2  ;
output wire [65:0] Final_58_F2_1_1  , Final_58_F2_1_2  , Final_58_F2_2_1  , Final_58_F2_2_2  ;
output wire [65:0] Final_58_F3_1_1  , Final_58_F3_1_2  , Final_58_F3_2_1  , Final_58_F3_2_2  ;
output wire [65:0] Final_58_F4_1_1  , Final_58_F4_1_2  , Final_58_F4_2_1  , Final_58_F4_2_2  ;
output wire [65:0] Final_59_F1_1_1  , Final_59_F1_1_2  , Final_59_F1_2_1  , Final_59_F1_2_2  ;
output wire [65:0] Final_59_F2_1_1  , Final_59_F2_1_2  , Final_59_F2_2_1  , Final_59_F2_2_2  ;
output wire [65:0] Final_59_F3_1_1  , Final_59_F3_1_2  , Final_59_F3_2_1  , Final_59_F3_2_2  ;
output wire [65:0] Final_59_F4_1_1  , Final_59_F4_1_2  , Final_59_F4_2_1  , Final_59_F4_2_2  ;
output wire [65:0] Final_60_F1_1_1  , Final_60_F1_1_2  , Final_60_F1_2_1  , Final_60_F1_2_2  ;
output wire [65:0] Final_60_F2_1_1  , Final_60_F2_1_2  , Final_60_F2_2_1  , Final_60_F2_2_2  ;
output wire [65:0] Final_60_F3_1_1  , Final_60_F3_1_2  , Final_60_F3_2_1  , Final_60_F3_2_2  ;
output wire [65:0] Final_60_F4_1_1  , Final_60_F4_1_2  , Final_60_F4_2_1  , Final_60_F4_2_2  ;
output wire [65:0] Final_61_F1_1_1  , Final_61_F1_1_2  , Final_61_F1_2_1  , Final_61_F1_2_2  ;
output wire [65:0] Final_61_F2_1_1  , Final_61_F2_1_2  , Final_61_F2_2_1  , Final_61_F2_2_2  ;
output wire [65:0] Final_61_F3_1_1  , Final_61_F3_1_2  , Final_61_F3_2_1  , Final_61_F3_2_2  ;
output wire [65:0] Final_61_F4_1_1  , Final_61_F4_1_2  , Final_61_F4_2_1  , Final_61_F4_2_2  ;
output wire [65:0] Final_62_F1_1_1  , Final_62_F1_1_2  , Final_62_F1_2_1  , Final_62_F1_2_2  ;
output wire [65:0] Final_62_F2_1_1  , Final_62_F2_1_2  , Final_62_F2_2_1  , Final_62_F2_2_2  ;
output wire [65:0] Final_62_F3_1_1  , Final_62_F3_1_2  , Final_62_F3_2_1  , Final_62_F3_2_2  ;
output wire [65:0] Final_62_F4_1_1  , Final_62_F4_1_2  , Final_62_F4_2_1  , Final_62_F4_2_2  ;
output wire [65:0] Final_63_F1_1_1  , Final_63_F1_1_2  , Final_63_F1_2_1  , Final_63_F1_2_2  ;
output wire [65:0] Final_63_F2_1_1  , Final_63_F2_1_2  , Final_63_F2_2_1  , Final_63_F2_2_2  ;
output wire [65:0] Final_63_F3_1_1  , Final_63_F3_1_2  , Final_63_F3_2_1  , Final_63_F3_2_2  ;
output wire [65:0] Final_63_F4_1_1  , Final_63_F4_1_2  , Final_63_F4_2_1  , Final_63_F4_2_2  ;
output wire [65:0] Final_64_F1_1_1  , Final_64_F1_1_2  , Final_64_F1_2_1  , Final_64_F1_2_2  ;
output wire [65:0] Final_64_F2_1_1  , Final_64_F2_1_2  , Final_64_F2_2_1  , Final_64_F2_2_2  ;
output wire [65:0] Final_64_F3_1_1  , Final_64_F3_1_2  , Final_64_F3_2_1  , Final_64_F3_2_2  ;
output wire [65:0] Final_64_F4_1_1  , Final_64_F4_1_2  , Final_64_F4_2_1  , Final_64_F4_2_2  ;
output wire [65:0] Final_65_F1_1_1  , Final_65_F1_1_2  , Final_65_F1_2_1  , Final_65_F1_2_2  ;
output wire [65:0] Final_65_F2_1_1  , Final_65_F2_1_2  , Final_65_F2_2_1  , Final_65_F2_2_2  ;
output wire [65:0] Final_65_F3_1_1  , Final_65_F3_1_2  , Final_65_F3_2_1  , Final_65_F3_2_2  ;
output wire [65:0] Final_65_F4_1_1  , Final_65_F4_1_2  , Final_65_F4_2_1  , Final_65_F4_2_2  ;
output wire [65:0] Final_66_F1_1_1  , Final_66_F1_1_2  , Final_66_F1_2_1  , Final_66_F1_2_2  ;
output wire [65:0] Final_66_F2_1_1  , Final_66_F2_1_2  , Final_66_F2_2_1  , Final_66_F2_2_2  ;
output wire [65:0] Final_66_F3_1_1  , Final_66_F3_1_2  , Final_66_F3_2_1  , Final_66_F3_2_2  ;
output wire [65:0] Final_66_F4_1_1  , Final_66_F4_1_2  , Final_66_F4_2_1  , Final_66_F4_2_2  ;
output wire [65:0] Final_67_F1_1_1  , Final_67_F1_1_2  , Final_67_F1_2_1  , Final_67_F1_2_2  ;
output wire [65:0] Final_67_F2_1_1  , Final_67_F2_1_2  , Final_67_F2_2_1  , Final_67_F2_2_2  ;
output wire [65:0] Final_67_F3_1_1  , Final_67_F3_1_2  , Final_67_F3_2_1  , Final_67_F3_2_2  ;
output wire [65:0] Final_67_F4_1_1  , Final_67_F4_1_2  , Final_67_F4_2_1  , Final_67_F4_2_2  ;
output wire [65:0] Final_68_F1_1_1  , Final_68_F1_1_2  , Final_68_F1_2_1  , Final_68_F1_2_2  ;
output wire [65:0] Final_68_F2_1_1  , Final_68_F2_1_2  , Final_68_F2_2_1  , Final_68_F2_2_2  ;
output wire [65:0] Final_68_F3_1_1  , Final_68_F3_1_2  , Final_68_F3_2_1  , Final_68_F3_2_2  ;
output wire [65:0] Final_68_F4_1_1  , Final_68_F4_1_2  , Final_68_F4_2_1  , Final_68_F4_2_2  ;
output wire [65:0] Final_69_F1_1_1  , Final_69_F1_1_2  , Final_69_F1_2_1  , Final_69_F1_2_2  ;
output wire [65:0] Final_69_F2_1_1  , Final_69_F2_1_2  , Final_69_F2_2_1  , Final_69_F2_2_2  ;
output wire [65:0] Final_69_F3_1_1  , Final_69_F3_1_2  , Final_69_F3_2_1  , Final_69_F3_2_2  ;
output wire [65:0] Final_69_F4_1_1  , Final_69_F4_1_2  , Final_69_F4_2_1  , Final_69_F4_2_2  ;
output wire [65:0] Final_70_F1_1_1  , Final_70_F1_1_2  , Final_70_F1_2_1  , Final_70_F1_2_2  ;
output wire [65:0] Final_70_F2_1_1  , Final_70_F2_1_2  , Final_70_F2_2_1  , Final_70_F2_2_2  ;
output wire [65:0] Final_70_F3_1_1  , Final_70_F3_1_2  , Final_70_F3_2_1  , Final_70_F3_2_2  ;
output wire [65:0] Final_70_F4_1_1  , Final_70_F4_1_2  , Final_70_F4_2_1  , Final_70_F4_2_2  ;
output wire [65:0] Final_71_F1_1_1  , Final_71_F1_1_2  , Final_71_F1_2_1  , Final_71_F1_2_2  ;
output wire [65:0] Final_71_F2_1_1  , Final_71_F2_1_2  , Final_71_F2_2_1  , Final_71_F2_2_2  ;
output wire [65:0] Final_71_F3_1_1  , Final_71_F3_1_2  , Final_71_F3_2_1  , Final_71_F3_2_2  ;
output wire [65:0] Final_71_F4_1_1  , Final_71_F4_1_2  , Final_71_F4_2_1  , Final_71_F4_2_2  ;
output wire [65:0] Final_72_F1_1_1  , Final_72_F1_1_2  , Final_72_F1_2_1  , Final_72_F1_2_2  ;
output wire [65:0] Final_72_F2_1_1  , Final_72_F2_1_2  , Final_72_F2_2_1  , Final_72_F2_2_2  ;
output wire [65:0] Final_72_F3_1_1  , Final_72_F3_1_2  , Final_72_F3_2_1  , Final_72_F3_2_2  ;
output wire [65:0] Final_72_F4_1_1  , Final_72_F4_1_2  , Final_72_F4_2_1  , Final_72_F4_2_2  ;
output wire [65:0] Final_73_F1_1_1  , Final_73_F1_1_2  , Final_73_F1_2_1  , Final_73_F1_2_2  ;
output wire [65:0] Final_73_F2_1_1  , Final_73_F2_1_2  , Final_73_F2_2_1  , Final_73_F2_2_2  ;
output wire [65:0] Final_73_F3_1_1  , Final_73_F3_1_2  , Final_73_F3_2_1  , Final_73_F3_2_2  ;
output wire [65:0] Final_73_F4_1_1  , Final_73_F4_1_2  , Final_73_F4_2_1  , Final_73_F4_2_2  ;
output wire [65:0] Final_74_F1_1_1  , Final_74_F1_1_2  , Final_74_F1_2_1  , Final_74_F1_2_2  ;
output wire [65:0] Final_74_F2_1_1  , Final_74_F2_1_2  , Final_74_F2_2_1  , Final_74_F2_2_2  ;
output wire [65:0] Final_74_F3_1_1  , Final_74_F3_1_2  , Final_74_F3_2_1  , Final_74_F3_2_2  ;
output wire [65:0] Final_74_F4_1_1  , Final_74_F4_1_2  , Final_74_F4_2_1  , Final_74_F4_2_2  ;
output wire [65:0] Final_75_F1_1_1  , Final_75_F1_1_2  , Final_75_F1_2_1  , Final_75_F1_2_2  ;
output wire [65:0] Final_75_F2_1_1  , Final_75_F2_1_2  , Final_75_F2_2_1  , Final_75_F2_2_2  ;
output wire [65:0] Final_75_F3_1_1  , Final_75_F3_1_2  , Final_75_F3_2_1  , Final_75_F3_2_2  ;
output wire [65:0] Final_75_F4_1_1  , Final_75_F4_1_2  , Final_75_F4_2_1  , Final_75_F4_2_2  ;
output wire [65:0] Final_76_F1_1_1  , Final_76_F1_1_2  , Final_76_F1_2_1  , Final_76_F1_2_2  ;
output wire [65:0] Final_76_F2_1_1  , Final_76_F2_1_2  , Final_76_F2_2_1  , Final_76_F2_2_2  ;
output wire [65:0] Final_76_F3_1_1  , Final_76_F3_1_2  , Final_76_F3_2_1  , Final_76_F3_2_2  ;
output wire [65:0] Final_76_F4_1_1  , Final_76_F4_1_2  , Final_76_F4_2_1  , Final_76_F4_2_2  ;
output wire [65:0] Final_77_F1_1_1  , Final_77_F1_1_2  , Final_77_F1_2_1  , Final_77_F1_2_2  ;
output wire [65:0] Final_77_F2_1_1  , Final_77_F2_1_2  , Final_77_F2_2_1  , Final_77_F2_2_2  ;
output wire [65:0] Final_77_F3_1_1  , Final_77_F3_1_2  , Final_77_F3_2_1  , Final_77_F3_2_2  ;
output wire [65:0] Final_77_F4_1_1  , Final_77_F4_1_2  , Final_77_F4_2_1  , Final_77_F4_2_2  ;
output wire [65:0] Final_78_F1_1_1  , Final_78_F1_1_2  , Final_78_F1_2_1  , Final_78_F1_2_2  ;
output wire [65:0] Final_78_F2_1_1  , Final_78_F2_1_2  , Final_78_F2_2_1  , Final_78_F2_2_2  ;
output wire [65:0] Final_78_F3_1_1  , Final_78_F3_1_2  , Final_78_F3_2_1  , Final_78_F3_2_2  ;
output wire [65:0] Final_78_F4_1_1  , Final_78_F4_1_2  , Final_78_F4_2_1  , Final_78_F4_2_2  ;
output wire [65:0] Final_79_F1_1_1  , Final_79_F1_1_2  , Final_79_F1_2_1  , Final_79_F1_2_2  ;
output wire [65:0] Final_79_F2_1_1  , Final_79_F2_1_2  , Final_79_F2_2_1  , Final_79_F2_2_2  ;
output wire [65:0] Final_79_F3_1_1  , Final_79_F3_1_2  , Final_79_F3_2_1  , Final_79_F3_2_2  ;
output wire [65:0] Final_79_F4_1_1  , Final_79_F4_1_2  , Final_79_F4_2_1  , Final_79_F4_2_2  ;
output wire [65:0] Final_80_F1_1_1  , Final_80_F1_1_2  , Final_80_F1_2_1  , Final_80_F1_2_2  ;
output wire [65:0] Final_80_F2_1_1  , Final_80_F2_1_2  , Final_80_F2_2_1  , Final_80_F2_2_2  ;
output wire [65:0] Final_80_F3_1_1  , Final_80_F3_1_2  , Final_80_F3_2_1  , Final_80_F3_2_2  ;
output wire [65:0] Final_80_F4_1_1  , Final_80_F4_1_2  , Final_80_F4_2_1  , Final_80_F4_2_2  ;
output wire [65:0] Final_81_F1_1_1  , Final_81_F1_1_2  , Final_81_F1_2_1  , Final_81_F1_2_2  ;
output wire [65:0] Final_81_F2_1_1  , Final_81_F2_1_2  , Final_81_F2_2_1  , Final_81_F2_2_2  ;
output wire [65:0] Final_81_F3_1_1  , Final_81_F3_1_2  , Final_81_F3_2_1  , Final_81_F3_2_2  ;
output wire [65:0] Final_81_F4_1_1  , Final_81_F4_1_2  , Final_81_F4_2_1  , Final_81_F4_2_2  ;
output wire [65:0] Final_82_F1_1_1  , Final_82_F1_1_2  , Final_82_F1_2_1  , Final_82_F1_2_2  ;
output wire [65:0] Final_82_F2_1_1  , Final_82_F2_1_2  , Final_82_F2_2_1  , Final_82_F2_2_2  ;
output wire [65:0] Final_82_F3_1_1  , Final_82_F3_1_2  , Final_82_F3_2_1  , Final_82_F3_2_2  ;
output wire [65:0] Final_82_F4_1_1  , Final_82_F4_1_2  , Final_82_F4_2_1  , Final_82_F4_2_2  ;
output wire [65:0] Final_83_F1_1_1  , Final_83_F1_1_2  , Final_83_F1_2_1  , Final_83_F1_2_2  ;
output wire [65:0] Final_83_F2_1_1  , Final_83_F2_1_2  , Final_83_F2_2_1  , Final_83_F2_2_2  ;
output wire [65:0] Final_83_F3_1_1  , Final_83_F3_1_2  , Final_83_F3_2_1  , Final_83_F3_2_2  ;
output wire [65:0] Final_83_F4_1_1  , Final_83_F4_1_2  , Final_83_F4_2_1  , Final_83_F4_2_2  ;
output wire [65:0] Final_84_F1_1_1  , Final_84_F1_1_2  , Final_84_F1_2_1  , Final_84_F1_2_2  ;
output wire [65:0] Final_84_F2_1_1  , Final_84_F2_1_2  , Final_84_F2_2_1  , Final_84_F2_2_2  ;
output wire [65:0] Final_84_F3_1_1  , Final_84_F3_1_2  , Final_84_F3_2_1  , Final_84_F3_2_2  ;
output wire [65:0] Final_84_F4_1_1  , Final_84_F4_1_2  , Final_84_F4_2_1  , Final_84_F4_2_2  ;
output wire [65:0] Final_85_F1_1_1  , Final_85_F1_1_2  , Final_85_F1_2_1  , Final_85_F1_2_2  ;
output wire [65:0] Final_85_F2_1_1  , Final_85_F2_1_2  , Final_85_F2_2_1  , Final_85_F2_2_2  ;
output wire [65:0] Final_85_F3_1_1  , Final_85_F3_1_2  , Final_85_F3_2_1  , Final_85_F3_2_2  ;
output wire [65:0] Final_85_F4_1_1  , Final_85_F4_1_2  , Final_85_F4_2_1  , Final_85_F4_2_2  ;
output wire [65:0] Final_86_F1_1_1  , Final_86_F1_1_2  , Final_86_F1_2_1  , Final_86_F1_2_2  ;
output wire [65:0] Final_86_F2_1_1  , Final_86_F2_1_2  , Final_86_F2_2_1  , Final_86_F2_2_2  ;
output wire [65:0] Final_86_F3_1_1  , Final_86_F3_1_2  , Final_86_F3_2_1  , Final_86_F3_2_2  ;
output wire [65:0] Final_86_F4_1_1  , Final_86_F4_1_2  , Final_86_F4_2_1  , Final_86_F4_2_2  ;
output wire [65:0] Final_87_F1_1_1  , Final_87_F1_1_2  , Final_87_F1_2_1  , Final_87_F1_2_2  ;
output wire [65:0] Final_87_F2_1_1  , Final_87_F2_1_2  , Final_87_F2_2_1  , Final_87_F2_2_2  ;
output wire [65:0] Final_87_F3_1_1  , Final_87_F3_1_2  , Final_87_F3_2_1  , Final_87_F3_2_2  ;
output wire [65:0] Final_87_F4_1_1  , Final_87_F4_1_2  , Final_87_F4_2_1  , Final_87_F4_2_2  ;
output wire [65:0] Final_88_F1_1_1  , Final_88_F1_1_2  , Final_88_F1_2_1  , Final_88_F1_2_2  ;
output wire [65:0] Final_88_F2_1_1  , Final_88_F2_1_2  , Final_88_F2_2_1  , Final_88_F2_2_2  ;
output wire [65:0] Final_88_F3_1_1  , Final_88_F3_1_2  , Final_88_F3_2_1  , Final_88_F3_2_2  ;
output wire [65:0] Final_88_F4_1_1  , Final_88_F4_1_2  , Final_88_F4_2_1  , Final_88_F4_2_2  ;
output wire [65:0] Final_89_F1_1_1  , Final_89_F1_1_2  , Final_89_F1_2_1  , Final_89_F1_2_2  ;
output wire [65:0] Final_89_F2_1_1  , Final_89_F2_1_2  , Final_89_F2_2_1  , Final_89_F2_2_2  ;
output wire [65:0] Final_89_F3_1_1  , Final_89_F3_1_2  , Final_89_F3_2_1  , Final_89_F3_2_2  ;
output wire [65:0] Final_89_F4_1_1  , Final_89_F4_1_2  , Final_89_F4_2_1  , Final_89_F4_2_2  ;
output wire [65:0] Final_90_F1_1_1  , Final_90_F1_1_2  , Final_90_F1_2_1  , Final_90_F1_2_2  ;
output wire [65:0] Final_90_F2_1_1  , Final_90_F2_1_2  , Final_90_F2_2_1  , Final_90_F2_2_2  ;
output wire [65:0] Final_90_F3_1_1  , Final_90_F3_1_2  , Final_90_F3_2_1  , Final_90_F3_2_2  ;
output wire [65:0] Final_90_F4_1_1  , Final_90_F4_1_2  , Final_90_F4_2_1  , Final_90_F4_2_2  ;
output wire [65:0] Final_91_F1_1_1  , Final_91_F1_1_2  , Final_91_F1_2_1  , Final_91_F1_2_2  ;
output wire [65:0] Final_91_F2_1_1  , Final_91_F2_1_2  , Final_91_F2_2_1  , Final_91_F2_2_2  ;
output wire [65:0] Final_91_F3_1_1  , Final_91_F3_1_2  , Final_91_F3_2_1  , Final_91_F3_2_2  ;
output wire [65:0] Final_91_F4_1_1  , Final_91_F4_1_2  , Final_91_F4_2_1  , Final_91_F4_2_2  ;
output wire [65:0] Final_92_F1_1_1  , Final_92_F1_1_2  , Final_92_F1_2_1  , Final_92_F1_2_2  ;
output wire [65:0] Final_92_F2_1_1  , Final_92_F2_1_2  , Final_92_F2_2_1  , Final_92_F2_2_2  ;
output wire [65:0] Final_92_F3_1_1  , Final_92_F3_1_2  , Final_92_F3_2_1  , Final_92_F3_2_2  ;
output wire [65:0] Final_92_F4_1_1  , Final_92_F4_1_2  , Final_92_F4_2_1  , Final_92_F4_2_2  ;
output wire [65:0] Final_93_F1_1_1  , Final_93_F1_1_2  , Final_93_F1_2_1  , Final_93_F1_2_2  ;
output wire [65:0] Final_93_F2_1_1  , Final_93_F2_1_2  , Final_93_F2_2_1  , Final_93_F2_2_2  ;
output wire [65:0] Final_93_F3_1_1  , Final_93_F3_1_2  , Final_93_F3_2_1  , Final_93_F3_2_2  ;
output wire [65:0] Final_93_F4_1_1  , Final_93_F4_1_2  , Final_93_F4_2_1  , Final_93_F4_2_2  ;
output wire [65:0] Final_94_F1_1_1  , Final_94_F1_1_2  , Final_94_F1_2_1  , Final_94_F1_2_2  ;
output wire [65:0] Final_94_F2_1_1  , Final_94_F2_1_2  , Final_94_F2_2_1  , Final_94_F2_2_2  ;
output wire [65:0] Final_94_F3_1_1  , Final_94_F3_1_2  , Final_94_F3_2_1  , Final_94_F3_2_2  ;
output wire [65:0] Final_94_F4_1_1  , Final_94_F4_1_2  , Final_94_F4_2_1  , Final_94_F4_2_2  ;
output wire [65:0] Final_95_F1_1_1  , Final_95_F1_1_2  , Final_95_F1_2_1  , Final_95_F1_2_2  ;
output wire [65:0] Final_95_F2_1_1  , Final_95_F2_1_2  , Final_95_F2_2_1  , Final_95_F2_2_2  ;
output wire [65:0] Final_95_F3_1_1  , Final_95_F3_1_2  , Final_95_F3_2_1  , Final_95_F3_2_2  ;
output wire [65:0] Final_95_F4_1_1  , Final_95_F4_1_2  , Final_95_F4_2_1  , Final_95_F4_2_2  ;
output wire [65:0] Final_96_F1_1_1  , Final_96_F1_1_2  , Final_96_F1_2_1  , Final_96_F1_2_2  ;
output wire [65:0] Final_96_F2_1_1  , Final_96_F2_1_2  , Final_96_F2_2_1  , Final_96_F2_2_2  ;
output wire [65:0] Final_96_F3_1_1  , Final_96_F3_1_2  , Final_96_F3_2_1  , Final_96_F3_2_2  ;
output wire [65:0] Final_96_F4_1_1  , Final_96_F4_1_2  , Final_96_F4_2_1  , Final_96_F4_2_2  ;
output wire [65:0] Final_97_F1_1_1  , Final_97_F1_1_2  , Final_97_F1_2_1  , Final_97_F1_2_2  ;
output wire [65:0] Final_97_F2_1_1  , Final_97_F2_1_2  , Final_97_F2_2_1  , Final_97_F2_2_2  ;
output wire [65:0] Final_97_F3_1_1  , Final_97_F3_1_2  , Final_97_F3_2_1  , Final_97_F3_2_2  ;
output wire [65:0] Final_97_F4_1_1  , Final_97_F4_1_2  , Final_97_F4_2_1  , Final_97_F4_2_2  ;
output wire [65:0] Final_98_F1_1_1  , Final_98_F1_1_2  , Final_98_F1_2_1  , Final_98_F1_2_2  ;
output wire [65:0] Final_98_F2_1_1  , Final_98_F2_1_2  , Final_98_F2_2_1  , Final_98_F2_2_2  ;
output wire [65:0] Final_98_F3_1_1  , Final_98_F3_1_2  , Final_98_F3_2_1  , Final_98_F3_2_2  ;
output wire [65:0] Final_98_F4_1_1  , Final_98_F4_1_2  , Final_98_F4_2_1  , Final_98_F4_2_2  ;
output wire [65:0] Final_99_F1_1_1  , Final_99_F1_1_2  , Final_99_F1_2_1  , Final_99_F1_2_2  ;
output wire [65:0] Final_99_F2_1_1  , Final_99_F2_1_2  , Final_99_F2_2_1  , Final_99_F2_2_2  ;
output wire [65:0] Final_99_F3_1_1  , Final_99_F3_1_2  , Final_99_F3_2_1  , Final_99_F3_2_2  ;
output wire [65:0] Final_99_F4_1_1  , Final_99_F4_1_2  , Final_99_F4_2_1  , Final_99_F4_2_2  ;
output wire [65:0] Final_100_F1_1_1  , Final_100_F1_1_2  , Final_100_F1_2_1  , Final_100_F1_2_2  ;
output wire [65:0] Final_100_F2_1_1  , Final_100_F2_1_2  , Final_100_F2_2_1  , Final_100_F2_2_2  ;
output wire [65:0] Final_100_F3_1_1  , Final_100_F3_1_2  , Final_100_F3_2_1  , Final_100_F3_2_2  ;
output wire [65:0] Final_100_F4_1_1  , Final_100_F4_1_2  , Final_100_F4_2_1  , Final_100_F4_2_2  ;
output wire [65:0] Final_101_F1_1_1  , Final_101_F1_1_2  , Final_101_F1_2_1  , Final_101_F1_2_2  ;
output wire [65:0] Final_101_F2_1_1  , Final_101_F2_1_2  , Final_101_F2_2_1  , Final_101_F2_2_2  ;
output wire [65:0] Final_101_F3_1_1  , Final_101_F3_1_2  , Final_101_F3_2_1  , Final_101_F3_2_2  ;
output wire [65:0] Final_101_F4_1_1  , Final_101_F4_1_2  , Final_101_F4_2_1  , Final_101_F4_2_2  ;
output wire [65:0] Final_102_F1_1_1  , Final_102_F1_1_2  , Final_102_F1_2_1  , Final_102_F1_2_2  ;
output wire [65:0] Final_102_F2_1_1  , Final_102_F2_1_2  , Final_102_F2_2_1  , Final_102_F2_2_2  ;
output wire [65:0] Final_102_F3_1_1  , Final_102_F3_1_2  , Final_102_F3_2_1  , Final_102_F3_2_2  ;
output wire [65:0] Final_102_F4_1_1  , Final_102_F4_1_2  , Final_102_F4_2_1  , Final_102_F4_2_2  ;
output wire [65:0] Final_103_F1_1_1  , Final_103_F1_1_2  , Final_103_F1_2_1  , Final_103_F1_2_2  ;
output wire [65:0] Final_103_F2_1_1  , Final_103_F2_1_2  , Final_103_F2_2_1  , Final_103_F2_2_2  ;
output wire [65:0] Final_103_F3_1_1  , Final_103_F3_1_2  , Final_103_F3_2_1  , Final_103_F3_2_2  ;
output wire [65:0] Final_103_F4_1_1  , Final_103_F4_1_2  , Final_103_F4_2_1  , Final_103_F4_2_2  ;
output wire [65:0] Final_104_F1_1_1  , Final_104_F1_1_2  , Final_104_F1_2_1  , Final_104_F1_2_2  ;
output wire [65:0] Final_104_F2_1_1  , Final_104_F2_1_2  , Final_104_F2_2_1  , Final_104_F2_2_2  ;
output wire [65:0] Final_104_F3_1_1  , Final_104_F3_1_2  , Final_104_F3_2_1  , Final_104_F3_2_2  ;
output wire [65:0] Final_104_F4_1_1  , Final_104_F4_1_2  , Final_104_F4_2_1  , Final_104_F4_2_2  ;
output wire [65:0] Final_105_F1_1_1  , Final_105_F1_1_2  , Final_105_F1_2_1  , Final_105_F1_2_2  ;
output wire [65:0] Final_105_F2_1_1  , Final_105_F2_1_2  , Final_105_F2_2_1  , Final_105_F2_2_2  ;
output wire [65:0] Final_105_F3_1_1  , Final_105_F3_1_2  , Final_105_F3_2_1  , Final_105_F3_2_2  ;
output wire [65:0] Final_105_F4_1_1  , Final_105_F4_1_2  , Final_105_F4_2_1  , Final_105_F4_2_2  ;
output wire [65:0] Final_106_F1_1_1  , Final_106_F1_1_2  , Final_106_F1_2_1  , Final_106_F1_2_2  ;
output wire [65:0] Final_106_F2_1_1  , Final_106_F2_1_2  , Final_106_F2_2_1  , Final_106_F2_2_2  ;
output wire [65:0] Final_106_F3_1_1  , Final_106_F3_1_2  , Final_106_F3_2_1  , Final_106_F3_2_2  ;
output wire [65:0] Final_106_F4_1_1  , Final_106_F4_1_2  , Final_106_F4_2_1  , Final_106_F4_2_2  ;
output wire [65:0] Final_107_F1_1_1  , Final_107_F1_1_2  , Final_107_F1_2_1  , Final_107_F1_2_2  ;
output wire [65:0] Final_107_F2_1_1  , Final_107_F2_1_2  , Final_107_F2_2_1  , Final_107_F2_2_2  ;
output wire [65:0] Final_107_F3_1_1  , Final_107_F3_1_2  , Final_107_F3_2_1  , Final_107_F3_2_2  ;
output wire [65:0] Final_107_F4_1_1  , Final_107_F4_1_2  , Final_107_F4_2_1  , Final_107_F4_2_2  ;
output wire [65:0] Final_108_F1_1_1  , Final_108_F1_1_2  , Final_108_F1_2_1  , Final_108_F1_2_2  ;
output wire [65:0] Final_108_F2_1_1  , Final_108_F2_1_2  , Final_108_F2_2_1  , Final_108_F2_2_2  ;
output wire [65:0] Final_108_F3_1_1  , Final_108_F3_1_2  , Final_108_F3_2_1  , Final_108_F3_2_2  ;
output wire [65:0] Final_108_F4_1_1  , Final_108_F4_1_2  , Final_108_F4_2_1  , Final_108_F4_2_2  ;
output wire [65:0] Final_109_F1_1_1  , Final_109_F1_1_2  , Final_109_F1_2_1  , Final_109_F1_2_2  ;
output wire [65:0] Final_109_F2_1_1  , Final_109_F2_1_2  , Final_109_F2_2_1  , Final_109_F2_2_2  ;
output wire [65:0] Final_109_F3_1_1  , Final_109_F3_1_2  , Final_109_F3_2_1  , Final_109_F3_2_2  ;
output wire [65:0] Final_109_F4_1_1  , Final_109_F4_1_2  , Final_109_F4_2_1  , Final_109_F4_2_2  ;
output wire [65:0] Final_110_F1_1_1  , Final_110_F1_1_2  , Final_110_F1_2_1  , Final_110_F1_2_2  ;
output wire [65:0] Final_110_F2_1_1  , Final_110_F2_1_2  , Final_110_F2_2_1  , Final_110_F2_2_2  ;
output wire [65:0] Final_110_F3_1_1  , Final_110_F3_1_2  , Final_110_F3_2_1  , Final_110_F3_2_2  ;
output wire [65:0] Final_110_F4_1_1  , Final_110_F4_1_2  , Final_110_F4_2_1  , Final_110_F4_2_2  ;
output wire [65:0] Final_111_F1_1_1  , Final_111_F1_1_2  , Final_111_F1_2_1  , Final_111_F1_2_2  ;
output wire [65:0] Final_111_F2_1_1  , Final_111_F2_1_2  , Final_111_F2_2_1  , Final_111_F2_2_2  ;
output wire [65:0] Final_111_F3_1_1  , Final_111_F3_1_2  , Final_111_F3_2_1  , Final_111_F3_2_2  ;
output wire [65:0] Final_111_F4_1_1  , Final_111_F4_1_2  , Final_111_F4_2_1  , Final_111_F4_2_2  ;
output wire [65:0] Final_112_F1_1_1  , Final_112_F1_1_2  , Final_112_F1_2_1  , Final_112_F1_2_2  ;
output wire [65:0] Final_112_F2_1_1  , Final_112_F2_1_2  , Final_112_F2_2_1  , Final_112_F2_2_2  ;
output wire [65:0] Final_112_F3_1_1  , Final_112_F3_1_2  , Final_112_F3_2_1  , Final_112_F3_2_2  ;
output wire [65:0] Final_112_F4_1_1  , Final_112_F4_1_2  , Final_112_F4_2_1  , Final_112_F4_2_2  ;
output wire [65:0] Final_113_F1_1_1  , Final_113_F1_1_2  , Final_113_F1_2_1  , Final_113_F1_2_2  ;
output wire [65:0] Final_113_F2_1_1  , Final_113_F2_1_2  , Final_113_F2_2_1  , Final_113_F2_2_2  ;
output wire [65:0] Final_113_F3_1_1  , Final_113_F3_1_2  , Final_113_F3_2_1  , Final_113_F3_2_2  ;
output wire [65:0] Final_113_F4_1_1  , Final_113_F4_1_2  , Final_113_F4_2_1  , Final_113_F4_2_2  ;
output wire [65:0] Final_114_F1_1_1  , Final_114_F1_1_2  , Final_114_F1_2_1  , Final_114_F1_2_2  ;
output wire [65:0] Final_114_F2_1_1  , Final_114_F2_1_2  , Final_114_F2_2_1  , Final_114_F2_2_2  ;
output wire [65:0] Final_114_F3_1_1  , Final_114_F3_1_2  , Final_114_F3_2_1  , Final_114_F3_2_2  ;
output wire [65:0] Final_114_F4_1_1  , Final_114_F4_1_2  , Final_114_F4_2_1  , Final_114_F4_2_2  ;
output wire [65:0] Final_115_F1_1_1  , Final_115_F1_1_2  , Final_115_F1_2_1  , Final_115_F1_2_2  ;
output wire [65:0] Final_115_F2_1_1  , Final_115_F2_1_2  , Final_115_F2_2_1  , Final_115_F2_2_2  ;
output wire [65:0] Final_115_F3_1_1  , Final_115_F3_1_2  , Final_115_F3_2_1  , Final_115_F3_2_2  ;
output wire [65:0] Final_115_F4_1_1  , Final_115_F4_1_2  , Final_115_F4_2_1  , Final_115_F4_2_2  ;
output wire [65:0] Final_116_F1_1_1  , Final_116_F1_1_2  , Final_116_F1_2_1  , Final_116_F1_2_2  ;
output wire [65:0] Final_116_F2_1_1  , Final_116_F2_1_2  , Final_116_F2_2_1  , Final_116_F2_2_2  ;
output wire [65:0] Final_116_F3_1_1  , Final_116_F3_1_2  , Final_116_F3_2_1  , Final_116_F3_2_2  ;
output wire [65:0] Final_116_F4_1_1  , Final_116_F4_1_2  , Final_116_F4_2_1  , Final_116_F4_2_2  ;
output wire [65:0] Final_117_F1_1_1  , Final_117_F1_1_2  , Final_117_F1_2_1  , Final_117_F1_2_2  ;
output wire [65:0] Final_117_F2_1_1  , Final_117_F2_1_2  , Final_117_F2_2_1  , Final_117_F2_2_2  ;
output wire [65:0] Final_117_F3_1_1  , Final_117_F3_1_2  , Final_117_F3_2_1  , Final_117_F3_2_2  ;
output wire [65:0] Final_117_F4_1_1  , Final_117_F4_1_2  , Final_117_F4_2_1  , Final_117_F4_2_2  ;
output wire [65:0] Final_118_F1_1_1  , Final_118_F1_1_2  , Final_118_F1_2_1  , Final_118_F1_2_2  ;
output wire [65:0] Final_118_F2_1_1  , Final_118_F2_1_2  , Final_118_F2_2_1  , Final_118_F2_2_2  ;
output wire [65:0] Final_118_F3_1_1  , Final_118_F3_1_2  , Final_118_F3_2_1  , Final_118_F3_2_2  ;
output wire [65:0] Final_118_F4_1_1  , Final_118_F4_1_2  , Final_118_F4_2_1  , Final_118_F4_2_2  ;
output wire [65:0] Final_119_F1_1_1  , Final_119_F1_1_2  , Final_119_F1_2_1  , Final_119_F1_2_2  ;
output wire [65:0] Final_119_F2_1_1  , Final_119_F2_1_2  , Final_119_F2_2_1  , Final_119_F2_2_2  ;
output wire [65:0] Final_119_F3_1_1  , Final_119_F3_1_2  , Final_119_F3_2_1  , Final_119_F3_2_2  ;
output wire [65:0] Final_119_F4_1_1  , Final_119_F4_1_2  , Final_119_F4_2_1  , Final_119_F4_2_2  ;
output wire [65:0] Final_120_F1_1_1  , Final_120_F1_1_2  , Final_120_F1_2_1  , Final_120_F1_2_2  ;
output wire [65:0] Final_120_F2_1_1  , Final_120_F2_1_2  , Final_120_F2_2_1  , Final_120_F2_2_2  ;
output wire [65:0] Final_120_F3_1_1  , Final_120_F3_1_2  , Final_120_F3_2_1  , Final_120_F3_2_2  ;
output wire [65:0] Final_120_F4_1_1  , Final_120_F4_1_2  , Final_120_F4_2_1  , Final_120_F4_2_2  ;
output wire [65:0] Final_121_F1_1_1  , Final_121_F1_1_2  , Final_121_F1_2_1  , Final_121_F1_2_2  ;
output wire [65:0] Final_121_F2_1_1  , Final_121_F2_1_2  , Final_121_F2_2_1  , Final_121_F2_2_2  ;
output wire [65:0] Final_121_F3_1_1  , Final_121_F3_1_2  , Final_121_F3_2_1  , Final_121_F3_2_2  ;
output wire [65:0] Final_121_F4_1_1  , Final_121_F4_1_2  , Final_121_F4_2_1  , Final_121_F4_2_2  ;
output wire [65:0] Final_122_F1_1_1  , Final_122_F1_1_2  , Final_122_F1_2_1  , Final_122_F1_2_2  ;
output wire [65:0] Final_122_F2_1_1  , Final_122_F2_1_2  , Final_122_F2_2_1  , Final_122_F2_2_2  ;
output wire [65:0] Final_122_F3_1_1  , Final_122_F3_1_2  , Final_122_F3_2_1  , Final_122_F3_2_2  ;
output wire [65:0] Final_122_F4_1_1  , Final_122_F4_1_2  , Final_122_F4_2_1  , Final_122_F4_2_2  ;
output wire [65:0] Final_123_F1_1_1  , Final_123_F1_1_2  , Final_123_F1_2_1  , Final_123_F1_2_2  ;
output wire [65:0] Final_123_F2_1_1  , Final_123_F2_1_2  , Final_123_F2_2_1  , Final_123_F2_2_2  ;
output wire [65:0] Final_123_F3_1_1  , Final_123_F3_1_2  , Final_123_F3_2_1  , Final_123_F3_2_2  ;
output wire [65:0] Final_123_F4_1_1  , Final_123_F4_1_2  , Final_123_F4_2_1  , Final_123_F4_2_2  ;
output wire [65:0] Final_124_F1_1_1  , Final_124_F1_1_2  , Final_124_F1_2_1  , Final_124_F1_2_2  ;
output wire [65:0] Final_124_F2_1_1  , Final_124_F2_1_2  , Final_124_F2_2_1  , Final_124_F2_2_2  ;
output wire [65:0] Final_124_F3_1_1  , Final_124_F3_1_2  , Final_124_F3_2_1  , Final_124_F3_2_2  ;
output wire [65:0] Final_124_F4_1_1  , Final_124_F4_1_2  , Final_124_F4_2_1  , Final_124_F4_2_2  ;
output wire [65:0] Final_125_F1_1_1  , Final_125_F1_1_2  , Final_125_F1_2_1  , Final_125_F1_2_2  ;
output wire [65:0] Final_125_F2_1_1  , Final_125_F2_1_2  , Final_125_F2_2_1  , Final_125_F2_2_2  ;
output wire [65:0] Final_125_F3_1_1  , Final_125_F3_1_2  , Final_125_F3_2_1  , Final_125_F3_2_2  ;
output wire [65:0] Final_125_F4_1_1  , Final_125_F4_1_2  , Final_125_F4_2_1  , Final_125_F4_2_2  ;
output wire [65:0] Final_126_F1_1_1  , Final_126_F1_1_2  , Final_126_F1_2_1  , Final_126_F1_2_2  ;
output wire [65:0] Final_126_F2_1_1  , Final_126_F2_1_2  , Final_126_F2_2_1  , Final_126_F2_2_2  ;
output wire [65:0] Final_126_F3_1_1  , Final_126_F3_1_2  , Final_126_F3_2_1  , Final_126_F3_2_2  ;
output wire [65:0] Final_126_F4_1_1  , Final_126_F4_1_2  , Final_126_F4_2_1  , Final_126_F4_2_2  ;
output wire [65:0] Final_127_F1_1_1  , Final_127_F1_1_2  , Final_127_F1_2_1  , Final_127_F1_2_2  ;
output wire [65:0] Final_127_F2_1_1  , Final_127_F2_1_2  , Final_127_F2_2_1  , Final_127_F2_2_2  ;
output wire [65:0] Final_127_F3_1_1  , Final_127_F3_1_2  , Final_127_F3_2_1  , Final_127_F3_2_2  ;
output wire [65:0] Final_127_F4_1_1  , Final_127_F4_1_2  , Final_127_F4_2_1  , Final_127_F4_2_2  ;
output wire [65:0] Final_128_F1_1_1  , Final_128_F1_1_2  , Final_128_F1_2_1  , Final_128_F1_2_2  ;
output wire [65:0] Final_128_F2_1_1  , Final_128_F2_1_2  , Final_128_F2_2_1  , Final_128_F2_2_2  ;
output wire [65:0] Final_128_F3_1_1  , Final_128_F3_1_2  , Final_128_F3_2_1  , Final_128_F3_2_2  ;
output wire [65:0] Final_128_F4_1_1  , Final_128_F4_1_2  , Final_128_F4_2_1  , Final_128_F4_2_2  ;
output wire [65:0] Final_129_F1_1_1  , Final_129_F1_1_2  , Final_129_F1_2_1  , Final_129_F1_2_2  ;
output wire [65:0] Final_129_F2_1_1  , Final_129_F2_1_2  , Final_129_F2_2_1  , Final_129_F2_2_2  ;
output wire [65:0] Final_129_F3_1_1  , Final_129_F3_1_2  , Final_129_F3_2_1  , Final_129_F3_2_2  ;
output wire [65:0] Final_129_F4_1_1  , Final_129_F4_1_2  , Final_129_F4_2_1  , Final_129_F4_2_2  ;
output wire [65:0] Final_130_F1_1_1  , Final_130_F1_1_2  , Final_130_F1_2_1  , Final_130_F1_2_2  ;
output wire [65:0] Final_130_F2_1_1  , Final_130_F2_1_2  , Final_130_F2_2_1  , Final_130_F2_2_2  ;
output wire [65:0] Final_130_F3_1_1  , Final_130_F3_1_2  , Final_130_F3_2_1  , Final_130_F3_2_2  ;
output wire [65:0] Final_130_F4_1_1  , Final_130_F4_1_2  , Final_130_F4_2_1  , Final_130_F4_2_2  ;
output wire [65:0] Final_131_F1_1_1  , Final_131_F1_1_2  , Final_131_F1_2_1  , Final_131_F1_2_2  ;
output wire [65:0] Final_131_F2_1_1  , Final_131_F2_1_2  , Final_131_F2_2_1  , Final_131_F2_2_2  ;
output wire [65:0] Final_131_F3_1_1  , Final_131_F3_1_2  , Final_131_F3_2_1  , Final_131_F3_2_2  ;
output wire [65:0] Final_131_F4_1_1  , Final_131_F4_1_2  , Final_131_F4_2_1  , Final_131_F4_2_2  ;
output wire [65:0] Final_132_F1_1_1  , Final_132_F1_1_2  , Final_132_F1_2_1  , Final_132_F1_2_2  ;
output wire [65:0] Final_132_F2_1_1  , Final_132_F2_1_2  , Final_132_F2_2_1  , Final_132_F2_2_2  ;
output wire [65:0] Final_132_F3_1_1  , Final_132_F3_1_2  , Final_132_F3_2_1  , Final_132_F3_2_2  ;
output wire [65:0] Final_132_F4_1_1  , Final_132_F4_1_2  , Final_132_F4_2_1  , Final_132_F4_2_2  ;
output wire [65:0] Final_133_F1_1_1  , Final_133_F1_1_2  , Final_133_F1_2_1  , Final_133_F1_2_2  ;
output wire [65:0] Final_133_F2_1_1  , Final_133_F2_1_2  , Final_133_F2_2_1  , Final_133_F2_2_2  ;
output wire [65:0] Final_133_F3_1_1  , Final_133_F3_1_2  , Final_133_F3_2_1  , Final_133_F3_2_2  ;
output wire [65:0] Final_133_F4_1_1  , Final_133_F4_1_2  , Final_133_F4_2_1  , Final_133_F4_2_2  ;
output wire [65:0] Final_134_F1_1_1  , Final_134_F1_1_2  , Final_134_F1_2_1  , Final_134_F1_2_2  ;
output wire [65:0] Final_134_F2_1_1  , Final_134_F2_1_2  , Final_134_F2_2_1  , Final_134_F2_2_2  ;
output wire [65:0] Final_134_F3_1_1  , Final_134_F3_1_2  , Final_134_F3_2_1  , Final_134_F3_2_2  ;
output wire [65:0] Final_134_F4_1_1  , Final_134_F4_1_2  , Final_134_F4_2_1  , Final_134_F4_2_2  ;
output wire [65:0] Final_135_F1_1_1  , Final_135_F1_1_2  , Final_135_F1_2_1  , Final_135_F1_2_2  ;
output wire [65:0] Final_135_F2_1_1  , Final_135_F2_1_2  , Final_135_F2_2_1  , Final_135_F2_2_2  ;
output wire [65:0] Final_135_F3_1_1  , Final_135_F3_1_2  , Final_135_F3_2_1  , Final_135_F3_2_2  ;
output wire [65:0] Final_135_F4_1_1  , Final_135_F4_1_2  , Final_135_F4_2_1  , Final_135_F4_2_2  ;
output wire [65:0] Final_136_F1_1_1  , Final_136_F1_1_2  , Final_136_F1_2_1  , Final_136_F1_2_2  ;
output wire [65:0] Final_136_F2_1_1  , Final_136_F2_1_2  , Final_136_F2_2_1  , Final_136_F2_2_2  ;
output wire [65:0] Final_136_F3_1_1  , Final_136_F3_1_2  , Final_136_F3_2_1  , Final_136_F3_2_2  ;
output wire [65:0] Final_136_F4_1_1  , Final_136_F4_1_2  , Final_136_F4_2_1  , Final_136_F4_2_2  ;
output wire [65:0] Final_137_F1_1_1  , Final_137_F1_1_2  , Final_137_F1_2_1  , Final_137_F1_2_2  ;
output wire [65:0] Final_137_F2_1_1  , Final_137_F2_1_2  , Final_137_F2_2_1  , Final_137_F2_2_2  ;
output wire [65:0] Final_137_F3_1_1  , Final_137_F3_1_2  , Final_137_F3_2_1  , Final_137_F3_2_2  ;
output wire [65:0] Final_137_F4_1_1  , Final_137_F4_1_2  , Final_137_F4_2_1  , Final_137_F4_2_2  ;
output wire [65:0] Final_138_F1_1_1  , Final_138_F1_1_2  , Final_138_F1_2_1  , Final_138_F1_2_2  ;
output wire [65:0] Final_138_F2_1_1  , Final_138_F2_1_2  , Final_138_F2_2_1  , Final_138_F2_2_2  ;
output wire [65:0] Final_138_F3_1_1  , Final_138_F3_1_2  , Final_138_F3_2_1  , Final_138_F3_2_2  ;
output wire [65:0] Final_138_F4_1_1  , Final_138_F4_1_2  , Final_138_F4_2_1  , Final_138_F4_2_2  ;
output wire [65:0] Final_139_F1_1_1  , Final_139_F1_1_2  , Final_139_F1_2_1  , Final_139_F1_2_2  ;
output wire [65:0] Final_139_F2_1_1  , Final_139_F2_1_2  , Final_139_F2_2_1  , Final_139_F2_2_2  ;
output wire [65:0] Final_139_F3_1_1  , Final_139_F3_1_2  , Final_139_F3_2_1  , Final_139_F3_2_2  ;
output wire [65:0] Final_139_F4_1_1  , Final_139_F4_1_2  , Final_139_F4_2_1  , Final_139_F4_2_2  ;
output wire [65:0] Final_140_F1_1_1  , Final_140_F1_1_2  , Final_140_F1_2_1  , Final_140_F1_2_2  ;
output wire [65:0] Final_140_F2_1_1  , Final_140_F2_1_2  , Final_140_F2_2_1  , Final_140_F2_2_2  ;
output wire [65:0] Final_140_F3_1_1  , Final_140_F3_1_2  , Final_140_F3_2_1  , Final_140_F3_2_2  ;
output wire [65:0] Final_140_F4_1_1  , Final_140_F4_1_2  , Final_140_F4_2_1  , Final_140_F4_2_2  ;
output wire [65:0] Final_141_F1_1_1  , Final_141_F1_1_2  , Final_141_F1_2_1  , Final_141_F1_2_2  ;
output wire [65:0] Final_141_F2_1_1  , Final_141_F2_1_2  , Final_141_F2_2_1  , Final_141_F2_2_2  ;
output wire [65:0] Final_141_F3_1_1  , Final_141_F3_1_2  , Final_141_F3_2_1  , Final_141_F3_2_2  ;
output wire [65:0] Final_141_F4_1_1  , Final_141_F4_1_2  , Final_141_F4_2_1  , Final_141_F4_2_2  ;
output wire [65:0] Final_142_F1_1_1  , Final_142_F1_1_2  , Final_142_F1_2_1  , Final_142_F1_2_2  ;
output wire [65:0] Final_142_F2_1_1  , Final_142_F2_1_2  , Final_142_F2_2_1  , Final_142_F2_2_2  ;
output wire [65:0] Final_142_F3_1_1  , Final_142_F3_1_2  , Final_142_F3_2_1  , Final_142_F3_2_2  ;
output wire [65:0] Final_142_F4_1_1  , Final_142_F4_1_2  , Final_142_F4_2_1  , Final_142_F4_2_2  ;
output wire [65:0] Final_143_F1_1_1  , Final_143_F1_1_2  , Final_143_F1_2_1  , Final_143_F1_2_2  ;
output wire [65:0] Final_143_F2_1_1  , Final_143_F2_1_2  , Final_143_F2_2_1  , Final_143_F2_2_2  ;
output wire [65:0] Final_143_F3_1_1  , Final_143_F3_1_2  , Final_143_F3_2_1  , Final_143_F3_2_2  ;
output wire [65:0] Final_143_F4_1_1  , Final_143_F4_1_2  , Final_143_F4_2_1  , Final_143_F4_2_2  ;
output wire [65:0] Final_144_F1_1_1  , Final_144_F1_1_2  , Final_144_F1_2_1  , Final_144_F1_2_2  ;
output wire [65:0] Final_144_F2_1_1  , Final_144_F2_1_2  , Final_144_F2_2_1  , Final_144_F2_2_2  ;
output wire [65:0] Final_144_F3_1_1  , Final_144_F3_1_2  , Final_144_F3_2_1  , Final_144_F3_2_2  ;
output wire [65:0] Final_144_F4_1_1  , Final_144_F4_1_2  , Final_144_F4_2_1  , Final_144_F4_2_2  ;


 */

//COUNTER_LAYER_6000_cycles count6000 (clk, bigaddress, Conv1LayerStart,tttt); 

COUNTER_LAYER_65536_cycles_NEW count65536 (clk, bigaddress, Conv1LayerStart, bigaddress340); //340 *144 = 48,960



wire rst;
//assign write2 = Conv1LayerFinish;
assign MAC_start = (counter >0) ?1'b1 :1'b0;//LayerStart;
assign MAC_end = (counter >338) ?1'b1 :1'b0;
assign rst = (counter ==9'b000000000)?1'b1 :1'b0; 

wire dummy;
reg resetTheCounter;


always @ (posedge clk)
begin
if (bigaddress ==   0) begin resetTheCounter <= 1; //340*0 = 0   bla_write<= 0;  BLA_address <= 0; 
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end

else if (bigaddress ==   340) begin resetTheCounter <= 1; //340*1 = 340
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   343) begin resetTheCounter <= 0;
write2_1  <= 1;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   680) begin resetTheCounter <= 1; //340*2 = 680
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   683) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 1;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   1020) begin resetTheCounter <= 1; //340*3 = 1020
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   1023) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 1;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   1360) begin resetTheCounter <= 1; //340*4 = 1360
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   1363) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 1;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   1700) begin resetTheCounter <= 1; //340*5 = 1700
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   1703) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 1;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   2040) begin resetTheCounter <= 1; //340*6 = 2040
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   2043) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 1;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   2380) begin resetTheCounter <= 1; //340*7 = 2380
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   2383) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 1;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   2720) begin resetTheCounter <= 1; //340*8 = 2720
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   2723) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 1;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   3060) begin resetTheCounter <= 1; //340*9 = 3060
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   3063) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 1;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   3400) begin resetTheCounter <= 1; //340*10 = 3400
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   3403) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 1;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   3740) begin resetTheCounter <= 1; //340*11 = 3740
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   3743) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 1;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   4080) begin resetTheCounter <= 1; //340*12 = 4080
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   4083) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 1;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   4420) begin resetTheCounter <= 1; //340*13 = 4420
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   4423) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 1;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   4760) begin resetTheCounter <= 1; //340*14 = 4760
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   4763) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 1;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   5100) begin resetTheCounter <= 1; //340*15 = 5100
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   5103) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 1;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   5440) begin resetTheCounter <= 1; //340*16 = 5440
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   5443) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 1;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   5780) begin resetTheCounter <= 1; //340*17 = 5780
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   5783) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 1;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   6120) begin resetTheCounter <= 1; //340*18 = 6120
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   6123) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 1;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   6460) begin resetTheCounter <= 1; //340*19 = 6460
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   6463) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 1;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   6800) begin resetTheCounter <= 1; //340*20 = 6800
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   6803) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 1;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   7140) begin resetTheCounter <= 1; //340*21 = 7140
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   7143) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 1;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   7480) begin resetTheCounter <= 1; //340*22 = 7480
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   7483) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 1;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   7820) begin resetTheCounter <= 1; //340*23 = 7820
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   7823) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 1;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   8160) begin resetTheCounter <= 1; //340*24 = 8160
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   8163) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 1;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   8500) begin resetTheCounter <= 1; //340*25 = 8500
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   8503) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 1;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   8840) begin resetTheCounter <= 1; //340*26 = 8840
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   8843) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 1;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   9180) begin resetTheCounter <= 1; //340*27 = 9180
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   9183) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 1;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   9520) begin resetTheCounter <= 1; //340*28 = 9520
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   9523) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 1;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   9860) begin resetTheCounter <= 1; //340*29 = 9860
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   9863) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 1;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   10200) begin resetTheCounter <= 1; //340*30 = 10200
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end

else if (bigaddress ==   10203) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 1;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   10540) begin resetTheCounter <= 1; //340*31 = 10540
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
///



else if (bigaddress ==   10543) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 1;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   10880) begin resetTheCounter <= 1; //340*32 = 10880
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   10883) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 1;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   11220) begin resetTheCounter <= 1; //340*33 = 11220
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   11223) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 1;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   11560) begin resetTheCounter <= 1; //340*34 = 11560
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   11563) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 1;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   11900) begin resetTheCounter <= 1; //340*35 = 11900
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   11903) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 1;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   12240) begin resetTheCounter <= 1; //340*36 = 12240
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   12243) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 1;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   12580) begin resetTheCounter <= 1; //340*37 = 12580
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   12583) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 1;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   12920) begin resetTheCounter <= 1; //340*38 = 12920
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   12923) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 1;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   13260) begin resetTheCounter <= 1; //340*39 = 13260
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   13263) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 1;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 

//40- 80

else if (bigaddress ==   13600) begin resetTheCounter <= 1; //340*40 = 13600
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   13603) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 1;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   13940) begin resetTheCounter <= 1; //340*41 = 13940
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   13943) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 1;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   14280) begin resetTheCounter <= 1; //340*42 = 14280
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   14283) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 1;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   14620) begin resetTheCounter <= 1; //340*43 = 14620
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   14623) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 1;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   14960) begin resetTheCounter <= 1; //340*44 = 14960
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   14963) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 1;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   15300) begin resetTheCounter <= 1; //340*45 = 15300
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   15303) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 1;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   15640) begin resetTheCounter <= 1; //340*46 = 15640
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   15643) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 1;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   15980) begin resetTheCounter <= 1; //340*47 = 15980
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   15983) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 1;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   16320) begin resetTheCounter <= 1; //340*48 = 16320
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   16323) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 1;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   16660) begin resetTheCounter <= 1; //340*49 = 16660
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   16663) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 1;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   17000) begin resetTheCounter <= 1; //340*50 = 17000
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   17003) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 1;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   17340) begin resetTheCounter <= 1; //340*51 = 17340
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   17343) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 1;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   17680) begin resetTheCounter <= 1; //340*52 = 17680
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   17683) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 1;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   18020) begin resetTheCounter <= 1; //340*53 = 18020
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   18023) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 1;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   18360) begin resetTheCounter <= 1; //340*54 = 18360
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   18363) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 1;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   18700) begin resetTheCounter <= 1; //340*55 = 18700
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   18703) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 1;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   19040) begin resetTheCounter <= 1; //340*56 = 19040
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   19043) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 1;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   19380) begin resetTheCounter <= 1; //340*57 = 19380
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   19383) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 1;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   19720) begin resetTheCounter <= 1; //340*58 = 19720
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   19723) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 1;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   20060) begin resetTheCounter <= 1; //340*59 = 20060
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   20063) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 1;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   20400) begin resetTheCounter <= 1; //340*60 = 20400
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   20403) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 1;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   20740) begin resetTheCounter <= 1; //340*61 = 20740
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   20743) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 1;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   21080) begin resetTheCounter <= 1; //340*62 = 21080
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   21083) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 1;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   21420) begin resetTheCounter <= 1; //340*63 = 21420
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   21423) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 1;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   21760) begin resetTheCounter <= 1; //340*64 = 21760
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   21763) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 1;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   22100) begin resetTheCounter <= 1; //340*65 = 22100
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   22103) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 1;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   22440) begin resetTheCounter <= 1; //340*66 = 22440
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   22443) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 1;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   22780) begin resetTheCounter <= 1; //340*67 = 22780
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   22783) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 1;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   23120) begin resetTheCounter <= 1; //340*68 = 23120
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   23123) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 1;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   23460) begin resetTheCounter <= 1; //340*69 = 23460
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   23463) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 1;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   23800) begin resetTheCounter <= 1; //340*70 = 23800
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   23803) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 1;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   24140) begin resetTheCounter <= 1; //340*71 = 24140
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   24143) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 1;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   24480) begin resetTheCounter <= 1; //340*72 = 24480
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   24483) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 1;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   24820) begin resetTheCounter <= 1; //340*73 = 24820
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   24823) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 1;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   25160) begin resetTheCounter <= 1; //340*74 = 25160
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   25163) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 1;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   25500) begin resetTheCounter <= 1; //340*75 = 25500
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   25503) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 1;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   25840) begin resetTheCounter <= 1; //340*76 = 25840
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   25843) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 1;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   26180) begin resetTheCounter <= 1; //340*77 = 26180
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   26183) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 1;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   26520) begin resetTheCounter <= 1; //340*78 = 26520
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   26523) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 1;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   26860) begin resetTheCounter <= 1; //340*79 = 26860
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   26863) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 1;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 

//80- 120


else if (bigaddress ==   27200) begin resetTheCounter <= 1; //340*80 = 27200
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   27203) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 1;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   27540) begin resetTheCounter <= 1; //340*81 = 27540
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   27543) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 1;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   27880) begin resetTheCounter <= 1; //340*82 = 27880
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   27883) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 1;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   28220) begin resetTheCounter <= 1; //340*83 = 28220
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   28223) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 1;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   28560) begin resetTheCounter <= 1; //340*84 = 28560
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   28563) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 1;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   28900) begin resetTheCounter <= 1; //340*85 = 28900
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   28903) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 1;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   29240) begin resetTheCounter <= 1; //340*86 = 29240
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   29243) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 1;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   29580) begin resetTheCounter <= 1; //340*87 = 29580
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   29583) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 1;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   29920) begin resetTheCounter <= 1; //340*88 = 29920
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   29923) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 1;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   30260) begin resetTheCounter <= 1; //340*89 = 30260
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   30263) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 1;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   30600) begin resetTheCounter <= 1; //340*90 = 30600
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   30603) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 1;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   30940) begin resetTheCounter <= 1; //340*91 = 30940
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   30943) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 1;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   31280) begin resetTheCounter <= 1; //340*92 = 31280
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   31283) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 1;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   31620) begin resetTheCounter <= 1; //340*93 = 31620
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   31623) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 1;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   31960) begin resetTheCounter <= 1; //340*94 = 31960
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   31963) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 1;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   32300) begin resetTheCounter <= 1; //340*95 = 32300
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   32303) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 1;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   32640) begin resetTheCounter <= 1; //340*96 = 32640
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   32643) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 1;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   32980) begin resetTheCounter <= 1; //340*97 = 32980
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   32983) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 1;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   33320) begin resetTheCounter <= 1; //340*98 = 33320
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   33323) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 1;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   33660) begin resetTheCounter <= 1; //340*99 = 33660
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   33663) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 1;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   34000) begin resetTheCounter <= 1; //340*100 = 34000
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   34003) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 1;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   34340) begin resetTheCounter <= 1; //340*101 = 34340
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   34343) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 1;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   34680) begin resetTheCounter <= 1; //340*102 = 34680
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   34683) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 1;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   35020) begin resetTheCounter <= 1; //340*103 = 35020
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   35023) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 1;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   35360) begin resetTheCounter <= 1; //340*104 = 35360
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   35363) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 1;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   35700) begin resetTheCounter <= 1; //340*105 = 35700
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   35703) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 1;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   36040) begin resetTheCounter <= 1; //340*106 = 36040
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   36043) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 1;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   36380) begin resetTheCounter <= 1; //340*107 = 36380
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   36383) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 1;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   36720) begin resetTheCounter <= 1; //340*108 = 36720
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   36723) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 1;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   37060) begin resetTheCounter <= 1; //340*109 = 37060
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   37063) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 1;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   37400) begin resetTheCounter <= 1; //340*110 = 37400
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   37403) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 1;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   37740) begin resetTheCounter <= 1; //340*111 = 37740
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   37743) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 1;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   38080) begin resetTheCounter <= 1; //340*112 = 38080
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   38083) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 1;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   38420) begin resetTheCounter <= 1; //340*113 = 38420
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   38423) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 1;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   38760) begin resetTheCounter <= 1; //340*114 = 38760
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   38763) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 1;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   39100) begin resetTheCounter <= 1; //340*115 = 39100
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   39103) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 1;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   39440) begin resetTheCounter <= 1; //340*116 = 39440
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   39443) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 1;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   39780) begin resetTheCounter <= 1; //340*117 = 39780
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   39783) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 1;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   40120) begin resetTheCounter <= 1; //340*118 = 40120
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   40123) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 1;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   40460) begin resetTheCounter <= 1; //340*119 = 40460
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   40463) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 1;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 

//120-144
else if (bigaddress ==   40800) begin resetTheCounter <= 1; //340*120 = 40800
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   40803) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 1;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   41140) begin resetTheCounter <= 1; //340*121 = 41140
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   41143) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 1;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   41480) begin resetTheCounter <= 1; //340*122 = 41480
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   41483) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 1;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   41820) begin resetTheCounter <= 1; //340*123 = 41820
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   41823) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 1;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   42160) begin resetTheCounter <= 1; //340*124 = 42160
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   42163) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 1;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   42500) begin resetTheCounter <= 1; //340*125 = 42500
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   42503) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 1;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   42840) begin resetTheCounter <= 1; //340*126 = 42840
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   42843) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 1;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   43180) begin resetTheCounter <= 1; //340*127 = 43180
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   43183) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 1;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   43520) begin resetTheCounter <= 1; //340*128 = 43520
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   43523) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 1;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   43860) begin resetTheCounter <= 1; //340*129 = 43860
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   43863) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 1;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   44200) begin resetTheCounter <= 1; //340*130 = 44200
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   44203) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 1;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   44540) begin resetTheCounter <= 1; //340*131 = 44540
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   44543) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 1;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   44880) begin resetTheCounter <= 1; //340*132 = 44880
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   44883) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 1;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   45220) begin resetTheCounter <= 1; //340*133 = 45220
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   45223) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 1;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   45560) begin resetTheCounter <= 1; //340*134 = 45560
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   45563) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 1;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   45900) begin resetTheCounter <= 1; //340*135 = 45900
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   45903) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 1;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   46240) begin resetTheCounter <= 1; //340*136 = 46240
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   46243) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 1;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   46580) begin resetTheCounter <= 1; //340*137 = 46580
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   46583) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 1;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   46920) begin resetTheCounter <= 1; //340*138 = 46920
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   46923) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 1;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   47260) begin resetTheCounter <= 1; //340*139 = 47260
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   47263) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 1;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   47600) begin resetTheCounter <= 1; //340*140 = 47600
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   47603) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 1;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   47940) begin resetTheCounter <= 1; //340*141 = 47940
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   47943) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 1;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   48280) begin resetTheCounter <= 1; //340*142 = 48280
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   48283) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 1;  write2_143  <= 0;  write2_144  <= 0; end
 
else if (bigaddress ==   48620) begin resetTheCounter <= 1; //340*143 = 48620
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   48623) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 1;  write2_144  <= 0; end
 
else if (bigaddress ==   48960) begin resetTheCounter <= 1; //340*144 = 48960
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
else if (bigaddress ==   48963) begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 1; end
 
else begin resetTheCounter <= 0;
write2_1  <= 0;  write2_2  <= 0;  write2_3  <= 0;  write2_4  <= 0;  write2_5  <= 0;  write2_6  <= 0;
write2_7  <= 0;  write2_8  <= 0;  write2_9  <= 0;  write2_10  <= 0;  write2_11  <= 0;  write2_12  <= 0;
write2_13  <= 0;  write2_14  <= 0;  write2_15  <= 0;  write2_16  <= 0;  write2_17  <= 0;  write2_18  <= 0;
write2_19  <= 0;  write2_20  <= 0;  write2_21  <= 0;  write2_22  <= 0;  write2_23  <= 0;  write2_24  <= 0;
write2_25  <= 0;  write2_26  <= 0;  write2_27  <= 0;  write2_28  <= 0;  write2_29  <= 0;  write2_30  <= 0;
write2_31  <= 0;  write2_32  <= 0;  write2_33  <= 0;  write2_34  <= 0;  write2_35  <= 0;  write2_36  <= 0;
write2_37  <= 0;  write2_38  <= 0;  write2_39  <= 0;  write2_40  <= 0;  write2_41  <= 0;  write2_42  <= 0;
write2_43  <= 0;  write2_44  <= 0;  write2_45  <= 0;  write2_46  <= 0;  write2_47  <= 0;  write2_48  <= 0;
write2_49  <= 0;  write2_50  <= 0;  write2_51  <= 0;  write2_52  <= 0;  write2_53  <= 0;  write2_54  <= 0;
write2_55  <= 0;  write2_56  <= 0;  write2_57  <= 0;  write2_58  <= 0;  write2_59  <= 0;  write2_60  <= 0;
write2_61  <= 0;  write2_62  <= 0;  write2_63  <= 0;  write2_64  <= 0;  write2_65  <= 0;  write2_66  <= 0;
write2_67  <= 0;  write2_68  <= 0;  write2_69  <= 0;  write2_70  <= 0;  write2_71  <= 0;  write2_72  <= 0;
write2_73  <= 0;  write2_74  <= 0;  write2_75  <= 0;  write2_76  <= 0;  write2_77  <= 0;  write2_78  <= 0;
write2_79  <= 0;  write2_80  <= 0;  write2_81  <= 0;  write2_82  <= 0;  write2_83  <= 0;  write2_84  <= 0;
write2_85  <= 0;  write2_86  <= 0;  write2_87  <= 0;  write2_88  <= 0;  write2_89  <= 0;  write2_90  <= 0;
write2_91  <= 0;  write2_92  <= 0;  write2_93  <= 0;  write2_94  <= 0;  write2_95  <= 0;  write2_96  <= 0;
write2_97  <= 0;  write2_98  <= 0;  write2_99  <= 0;  write2_100  <= 0;  write2_101  <= 0;  write2_102  <= 0;
write2_103  <= 0;  write2_104  <= 0;  write2_105  <= 0;  write2_106  <= 0;  write2_107  <= 0;  write2_108  <= 0;
write2_109  <= 0;  write2_110  <= 0;  write2_111  <= 0;  write2_112  <= 0;  write2_113  <= 0;  write2_114  <= 0;
write2_115  <= 0;  write2_116  <= 0;  write2_117  <= 0;  write2_118  <= 0;  write2_119  <= 0;  write2_120  <= 0;
write2_121  <= 0;  write2_122  <= 0;  write2_123  <= 0;  write2_124  <= 0;  write2_125  <= 0;  write2_126  <= 0;
write2_127  <= 0;  write2_128  <= 0;  write2_129  <= 0;  write2_130  <= 0;  write2_131  <= 0;  write2_132  <= 0;
write2_133  <= 0;  write2_134  <= 0;  write2_135  <= 0;  write2_136  <= 0;  write2_137  <= 0;  write2_138  <= 0;
write2_139  <= 0;  write2_140  <= 0;  write2_141  <= 0;  write2_142  <= 0;  write2_143  <= 0;  write2_144  <= 0; end
 
end



//assign Conv1LayerFinish = (bigaddress == 48962) ?1'b1 :1'b0;
assign MAX1LayerFinish = (bigaddress == 48962) ?1'b1 :1'b0;

COUNTER_LAYER_340_cycles Counter340 (clk, resetTheCounter, counter, Conv1LayerStart ,dummy);
//resetTheCounter
ROM_26x66bit_F1 FilterWeights1 (clk, counter, ROMout1 );
ROM_26x66bit_F2 FilterWeights2 (clk, counter, ROMout2 );
ROM_26x66bit_F3 FilterWeights3 (clk, counter, ROMout3 );
ROM_26x66bit_F4 FilterWeights4 (clk, counter, ROMout4 );


main_fsm_CONV ConvStateMachine (clk, rst, counter, address);



//36 16*26 mux

//26 * 16 * 1 = 416 * 1 (36 muxes from this) 
//we don't need all this enough 100 * 1 (36 muxes from this) 


WireDivision mux1_1_1_1(  DataOut0, DataOut2, DataOut4, DataOut6, DataOut8, DataOut10, DataOut12, DataOut14, DataOut16, DataOut18, DataOut20, DataOut22, DataOut56, DataOut58, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut112, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut168, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut224, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut280, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut336, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut392, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut448, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut504, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut560, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut616, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638,  bigaddress340, Super_1_1_1_1);
WireDivision mux1_2_1_1(  DataOut1, DataOut3, DataOut5, DataOut7, DataOut9, DataOut11, DataOut13, DataOut15, DataOut17, DataOut19, DataOut21, DataOut23, DataOut57, DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut113, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut169, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut225, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut281, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut337, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut393, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut449, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut505, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut561, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut617, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639,  bigaddress340, Super_1_2_1_1);
WireDivision mux1_3_1_1(  DataOut2, DataOut4, DataOut6, DataOut8, DataOut10, DataOut12, DataOut14, DataOut16, DataOut18, DataOut20, DataOut22, DataOut24, DataOut58, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640 , bigaddress340, Super_1_3_1_1);
WireDivision mux1_4_1_1(  DataOut3, DataOut5, DataOut7, DataOut9, DataOut11, DataOut13, DataOut15, DataOut17, DataOut19, DataOut21, DataOut23, DataOut25, DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut81, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641,  bigaddress340, Super_1_4_1_1);
WireDivision mux1_5_1_1(  DataOut4, DataOut6, DataOut8, DataOut10, DataOut12, DataOut14, DataOut16, DataOut18, DataOut20, DataOut22, DataOut24, DataOut26, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut82, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut138, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut194, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut250, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut306, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut362, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut418, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut474, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut530, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut586, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut642,  bigaddress340, Super_1_5_1_1);

WireDivision mux2_1_1_1(  DataOut28, DataOut30, DataOut32, DataOut34, DataOut36, DataOut38, DataOut40, DataOut42, DataOut44, DataOut46, DataOut48, DataOut50, DataOut84, DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut140, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut196, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut252, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut308, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut364, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut420, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut476, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut532, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut588, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut644, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666,  bigaddress340, Super_2_1_1_1);
WireDivision mux2_2_1_1(  DataOut29, DataOut31, DataOut33, DataOut35, DataOut37, DataOut39, DataOut41, DataOut43, DataOut45, DataOut47, DataOut49, DataOut51, DataOut85, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut141, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut197, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut253, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut309, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut365, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut421, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut477, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut533, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut589, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut645, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667,  bigaddress340, Super_2_2_1_1);
WireDivision mux2_3_1_1(  DataOut30, DataOut32, DataOut34, DataOut36, DataOut38, DataOut40, DataOut42, DataOut44, DataOut46, DataOut48, DataOut50, DataOut52, DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668,  bigaddress340, Super_2_3_1_1);
WireDivision mux2_4_1_1(  DataOut31, DataOut33, DataOut35, DataOut37, DataOut39, DataOut41, DataOut43, DataOut45, DataOut47, DataOut49, DataOut51, DataOut53, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669,  bigaddress340, Super_2_4_1_1);
WireDivision mux2_5_1_1(  DataOut32, DataOut34, DataOut36, DataOut38, DataOut40, DataOut42, DataOut44, DataOut46, DataOut48, DataOut50, DataOut52, DataOut54, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut110, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670,  bigaddress340, Super_2_5_1_1);

WireDivision mux3_1_1_1(  DataOut56, DataOut58, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut112, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut168, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut224, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut280, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut336, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut392, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut448, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut504, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut560, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut616, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut672, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694,  bigaddress340, Super_3_1_1_1);
WireDivision mux3_2_1_1(  DataOut57, DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut113, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut169, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut225, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut281, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut337, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut393, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut449, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut505, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut561, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut617, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut673, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695,  bigaddress340, Super_3_2_1_1);
WireDivision mux3_3_1_1(  DataOut58, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696,  bigaddress340, Super_3_3_1_1);
WireDivision mux3_4_1_1(  DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut81, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697,  bigaddress340, Super_3_4_1_1);
WireDivision mux3_5_1_1(  DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut82, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut138, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut194, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut250, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut306, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut362, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut418, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut474, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut530, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut586, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut642, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut698,  bigaddress340, Super_3_5_1_1);

WireDivision mux4_1_1_1(  DataOut84, DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut140, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut196, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut252, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut308, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut364, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut420, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut476, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut532, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut588, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut644, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut700, DataOut702, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722,  bigaddress340, Super_4_1_1_1);
WireDivision mux4_2_1_1(  DataOut85, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut141, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut197, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut253, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut309, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut365, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut421, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut477, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut533, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut589, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut645, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut701, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723,  bigaddress340, Super_4_2_1_1);
WireDivision mux4_3_1_1(  DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut702, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724,  bigaddress340, Super_4_3_1_1);
WireDivision mux4_4_1_1(  DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725,  bigaddress340, Super_4_4_1_1);
WireDivision mux4_5_1_1(  DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut110, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724, DataOut726,  bigaddress340, Super_4_5_1_1);

WireDivision mux5_1_1_1(  DataOut112, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut168, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut224, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut280, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut336, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut392, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut448, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut504, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut560, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut616, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut672, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut728, DataOut730, DataOut732, DataOut734, DataOut736, DataOut738, DataOut740, DataOut742, DataOut744, DataOut746, DataOut748, DataOut750,  bigaddress340, Super_5_1_1_1);
WireDivision mux5_2_1_1(  DataOut113, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut169, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut225, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut281, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut337, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut393, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut449, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut505, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut561, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut617, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut673, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut729, DataOut731, DataOut733, DataOut735, DataOut737, DataOut739, DataOut741, DataOut743, DataOut745, DataOut747, DataOut749, DataOut751,  bigaddress340, Super_5_2_1_1);
WireDivision mux5_3_1_1(  DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut730, DataOut732, DataOut734, DataOut736, DataOut738, DataOut740, DataOut742, DataOut744, DataOut746, DataOut748, DataOut750, DataOut752,  bigaddress340, Super_5_3_1_1);
WireDivision mux5_4_1_1(  DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697, DataOut731, DataOut733, DataOut735, DataOut737, DataOut739, DataOut741, DataOut743, DataOut745, DataOut747, DataOut749, DataOut751, DataOut753,  bigaddress340, Super_5_4_1_1);
WireDivision mux5_5_1_1(  DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut138, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut194, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut250, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut306, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut362, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut418, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut474, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut530, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut586, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut642, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut698, DataOut732, DataOut734, DataOut736, DataOut738, DataOut740, DataOut742, DataOut744, DataOut746, DataOut748, DataOut750, DataOut752, DataOut754,  bigaddress340, Super_5_5_1_1);



WireDivision mux1_1_1_2(  DataOut1, DataOut3, DataOut5, DataOut7, DataOut9, DataOut11, DataOut13, DataOut15, DataOut17, DataOut19, DataOut21, DataOut23, DataOut57, DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut113, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut169, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut225, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut281, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut337, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut393, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut449, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut505, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut561, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut617, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639,  bigaddress340, Super_1_1_1_2);
WireDivision mux1_2_1_2(  DataOut2, DataOut4, DataOut6, DataOut8, DataOut10, DataOut12, DataOut14, DataOut16, DataOut18, DataOut20, DataOut22, DataOut24, DataOut58, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640,  bigaddress340, Super_1_2_1_2);
WireDivision mux1_3_1_2(  DataOut3, DataOut5, DataOut7, DataOut9, DataOut11, DataOut13, DataOut15, DataOut17, DataOut19, DataOut21, DataOut23, DataOut25, DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut81, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641,  bigaddress340, Super_1_3_1_2);
WireDivision mux1_4_1_2(  DataOut4, DataOut6, DataOut8, DataOut10, DataOut12, DataOut14, DataOut16, DataOut18, DataOut20, DataOut22, DataOut24, DataOut26, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut82, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut138, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut194, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut250, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut306, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut362, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut418, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut474, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut530, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut586, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut642,  bigaddress340, Super_1_4_1_2);
WireDivision mux1_5_1_2(  DataOut5, DataOut7, DataOut9, DataOut11, DataOut13, DataOut15, DataOut17, DataOut19, DataOut21, DataOut23, DataOut25, DataOut27, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut81, DataOut83, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut139, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut195, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut251, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut307, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut363, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut419, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut475, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut531, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut587, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut643,  bigaddress340, Super_1_5_1_2);


WireDivision mux2_1_1_2(  DataOut29, DataOut31, DataOut33, DataOut35, DataOut37, DataOut39, DataOut41, DataOut43, DataOut45, DataOut47, DataOut49, DataOut51, DataOut85, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut141, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut197, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut253, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut309, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut365, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut421, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut477, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut533, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut589, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut645, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667,  bigaddress340, Super_2_1_1_2);
WireDivision mux2_2_1_2(  DataOut30, DataOut32, DataOut34, DataOut36, DataOut38, DataOut40, DataOut42, DataOut44, DataOut46, DataOut48, DataOut50, DataOut52, DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668,  bigaddress340, Super_2_2_1_2);
WireDivision mux2_3_1_2(  DataOut31, DataOut33, DataOut35, DataOut37, DataOut39, DataOut41, DataOut43, DataOut45, DataOut47, DataOut49, DataOut51, DataOut53, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, bigaddress340, Super_2_3_1_2);
WireDivision mux2_4_1_2(  DataOut32, DataOut34, DataOut36, DataOut38, DataOut40, DataOut42, DataOut44, DataOut46, DataOut48, DataOut50, DataOut52, DataOut54, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut110, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670, bigaddress340, Super_2_4_1_2);
WireDivision mux2_5_1_2(  DataOut33, DataOut35, DataOut37, DataOut39, DataOut41, DataOut43, DataOut45, DataOut47, DataOut49, DataOut51, DataOut53, DataOut55, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut111, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut167, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut223, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut279, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut335, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut391, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut447, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut503, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut559, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut615, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut671, bigaddress340, Super_2_5_1_2);

WireDivision mux3_1_1_2(  DataOut57, DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut113, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut169, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut225, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut281, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut337, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut393, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut449, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut505, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut561, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut617, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut673, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695,  bigaddress340, Super_3_1_1_2);
WireDivision mux3_2_1_2(  DataOut58, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696,  bigaddress340, Super_3_2_1_2);
WireDivision mux3_3_1_2(  DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut81, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697,  bigaddress340, Super_3_3_1_2);
WireDivision mux3_4_1_2(  DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut82, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut138, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut194, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut250, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut306, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut362, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut418, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut474, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut530, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut586, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut642, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut698,  bigaddress340, Super_3_4_1_2);
WireDivision mux3_5_1_2(  DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut81, DataOut83, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut139, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut195, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut251, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut307, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut363, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut419, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut475, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut531, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut587, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut643, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697, DataOut699,  bigaddress340, Super_3_5_1_2);

WireDivision mux4_1_1_2( DataOut85, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut141, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut197, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut253, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut309, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut365, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut421, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut477, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut533, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut589, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut645, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut701, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723,   bigaddress340, Super_4_1_1_2);
WireDivision mux4_2_1_2( DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut702, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724,   bigaddress340, Super_4_2_1_2);
WireDivision mux4_3_1_2( DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725,   bigaddress340, Super_4_3_1_2);
WireDivision mux4_4_1_2( DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut110, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724, DataOut726,   bigaddress340, Super_4_4_1_2);
WireDivision mux4_5_1_2( DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut111, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut167, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut223, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut279, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut335, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut391, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut447, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut503, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut559, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut615, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut671, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725, DataOut727,   bigaddress340, Super_4_5_1_2);

WireDivision mux5_1_1_2(  DataOut113, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut169, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut225, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut281, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut337, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut393, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut449, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut505, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut561, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut617, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut673, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut729, DataOut731, DataOut733, DataOut735, DataOut737, DataOut739, DataOut741, DataOut743, DataOut745, DataOut747, DataOut749, DataOut751,  bigaddress340, Super_5_1_1_2);
WireDivision mux5_2_1_2(  DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut730, DataOut732, DataOut734, DataOut736, DataOut738, DataOut740, DataOut742, DataOut744, DataOut746, DataOut748, DataOut750, DataOut752,  bigaddress340, Super_5_2_1_2);
WireDivision mux5_3_1_2( DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697, DataOut731, DataOut733, DataOut735, DataOut737, DataOut739, DataOut741, DataOut743, DataOut745, DataOut747, DataOut749, DataOut751, DataOut753,   bigaddress340, Super_5_3_1_2);
WireDivision mux5_4_1_2(  DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut138, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut194, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut250, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut306, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut362, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut418, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut474, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut530, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut586, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut642, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut698, DataOut732, DataOut734, DataOut736, DataOut738, DataOut740, DataOut742, DataOut744, DataOut746, DataOut748, DataOut750, DataOut752, DataOut754,  bigaddress340, Super_5_4_1_2);
WireDivision mux5_5_1_2(  DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut139, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut195, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut251, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut307, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut363, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut419, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut475, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut531, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut587, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut643, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697, DataOut699, DataOut733, DataOut735, DataOut737, DataOut739, DataOut741, DataOut743, DataOut745, DataOut747, DataOut749, DataOut751, DataOut753, DataOut755,  bigaddress340, Super_5_5_1_2);



WireDivision mux1_1_2_1(  DataOut28, DataOut30, DataOut32, DataOut34, DataOut36, DataOut38, DataOut40, DataOut42, DataOut44, DataOut46, DataOut48, DataOut50, DataOut84, DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut140, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut196, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut252, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut308, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut364, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut420, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut476, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut532, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut588, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut644, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666,  bigaddress340, Super_1_1_2_1);
WireDivision mux1_2_2_1(  DataOut29, DataOut31, DataOut33, DataOut35, DataOut37, DataOut39, DataOut41, DataOut43, DataOut45, DataOut47, DataOut49, DataOut51, DataOut85, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut141, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut197, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut253, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut309, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut365, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut421, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut477, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut533, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut589, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut645, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667,  bigaddress340, Super_1_2_2_1);
WireDivision mux1_3_2_1(  DataOut30, DataOut32, DataOut34, DataOut36, DataOut38, DataOut40, DataOut42, DataOut44, DataOut46, DataOut48, DataOut50, DataOut52, DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668,  bigaddress340, Super_1_3_2_1);
WireDivision mux1_4_2_1(  DataOut31, DataOut33, DataOut35, DataOut37, DataOut39, DataOut41, DataOut43, DataOut45, DataOut47, DataOut49, DataOut51, DataOut53, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669,  bigaddress340, Super_1_4_2_1);
WireDivision mux1_5_2_1(  DataOut32, DataOut34, DataOut36, DataOut38, DataOut40, DataOut42, DataOut44, DataOut46, DataOut48, DataOut50, DataOut52, DataOut54, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut110, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670,  bigaddress340, Super_1_5_2_1);

WireDivision mux2_1_2_1(  DataOut56, DataOut58, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut112, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut168, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut224, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut280, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut336, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut392, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut448, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut504, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut560, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut616, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut672, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, bigaddress340, Super_2_1_2_1);
WireDivision mux2_2_2_1(  DataOut57, DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut113, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut169, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut225, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut281, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut337, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut393, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut449, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut505, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut561, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut617, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut673, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695,  bigaddress340, Super_2_2_2_1);
WireDivision mux2_3_2_1(  DataOut58, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696,  bigaddress340, Super_2_3_2_1);
WireDivision mux2_4_2_1(  DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut81, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697,  bigaddress340, Super_2_4_2_1);
WireDivision mux2_5_2_1(  DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut82, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut138, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut194, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut250, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut306, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut362, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut418, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut474, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut530, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut586, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut642, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut698,  bigaddress340, Super_2_5_2_1);

WireDivision mux3_1_2_1( DataOut84, DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut140, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut196, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut252, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut308, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut364, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut420, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut476, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut532, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut588, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut644, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut700, DataOut702, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, bigaddress340, Super_3_1_2_1);
WireDivision mux3_2_2_1( DataOut85, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut141, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut197, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut253, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut309, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut365, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut421, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut477, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut533, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut589, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut645, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut701, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, bigaddress340, Super_3_2_2_1);
WireDivision mux3_3_2_1( DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut702, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724,   bigaddress340, Super_3_3_2_1);
WireDivision mux3_4_2_1( DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725, bigaddress340, Super_3_4_2_1); // DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725,   bigaddress340, Super_3_4_2_1);
WireDivision mux3_5_2_1( DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut110, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724, DataOut726,bigaddress340, Super_3_5_2_1);// DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut110, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724, DataOut726,   bigaddress340, Super_3_5_2_1);

WireDivision mux4_1_2_1( DataOut112, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut168, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut224, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut280, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut336, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut392, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut448, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut504, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut560, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut616, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut672, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut728, DataOut730, DataOut732, DataOut734, DataOut736, DataOut738, DataOut740, DataOut742, DataOut744, DataOut746, DataOut748, DataOut750,   bigaddress340, Super_4_1_2_1);
WireDivision mux4_2_2_1( DataOut113, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut169, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut225, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut281, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut337, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut393, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut449, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut505, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut561, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut617, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut673, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut729, DataOut731, DataOut733, DataOut735, DataOut737, DataOut739, DataOut741, DataOut743, DataOut745, DataOut747, DataOut749, DataOut751,   bigaddress340, Super_4_2_2_1);
WireDivision mux4_3_2_1( DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut730, DataOut732, DataOut734, DataOut736, DataOut738, DataOut740, DataOut742, DataOut744, DataOut746, DataOut748, DataOut750, DataOut752,   bigaddress340, Super_4_3_2_1);
WireDivision mux4_4_2_1( DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697, DataOut731, DataOut733, DataOut735, DataOut737, DataOut739, DataOut741, DataOut743, DataOut745, DataOut747, DataOut749, DataOut751, DataOut753,   bigaddress340, Super_4_4_2_1);
WireDivision mux4_5_2_1( DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut138, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut194, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut250, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut306, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut362, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut418, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut474, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut530, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut586, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut642, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut698, DataOut732, DataOut734, DataOut736, DataOut738, DataOut740, DataOut742, DataOut744, DataOut746, DataOut748, DataOut750, DataOut752, DataOut754,   bigaddress340, Super_4_5_2_1);

WireDivision mux5_1_2_1(  DataOut140, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut196, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut252, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut308, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut364, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut420, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut476, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut532, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut588, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut644, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut700, DataOut702, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut756, DataOut758, DataOut760, DataOut762, DataOut764, DataOut766, DataOut768, DataOut770, DataOut772, DataOut774, DataOut776, DataOut778,  bigaddress340, Super_5_1_2_1);
WireDivision mux5_2_2_1(  DataOut141, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut197, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut253, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut309, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut365, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut421, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut477, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut533, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut589, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut645, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut701, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut757, DataOut759, DataOut761, DataOut763, DataOut765, DataOut767, DataOut769, DataOut771, DataOut773, DataOut775, DataOut777, DataOut779,  bigaddress340, Super_5_2_2_1);
WireDivision mux5_3_2_1(  DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut702, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724, DataOut758, DataOut760, DataOut762, DataOut764, DataOut766, DataOut768, DataOut770, DataOut772, DataOut774, DataOut776, DataOut778, DataOut780,  bigaddress340, Super_5_3_2_1);
WireDivision mux5_4_2_1(  DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725, DataOut759, DataOut761, DataOut763, DataOut765, DataOut767, DataOut769, DataOut771, DataOut773, DataOut775, DataOut777, DataOut779, DataOut781,  bigaddress340, Super_5_4_2_1);
WireDivision mux5_5_2_1(  DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724, DataOut726, DataOut760, DataOut762, DataOut764, DataOut766, DataOut768, DataOut770, DataOut772, DataOut774, DataOut776, DataOut778, DataOut780, DataOut782,  bigaddress340, Super_5_5_2_1);



WireDivision mux1_1_2_2(  DataOut29, DataOut31, DataOut33, DataOut35, DataOut37, DataOut39, DataOut41, DataOut43, DataOut45, DataOut47, DataOut49, DataOut51, DataOut85, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut141, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut197, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut253, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut309, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut365, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut421, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut477, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut533, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut589, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut645, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667,  bigaddress340, Super_1_1_2_2);
WireDivision mux1_2_2_2(  DataOut30, DataOut32, DataOut34, DataOut36, DataOut38, DataOut40, DataOut42, DataOut44, DataOut46, DataOut48, DataOut50, DataOut52, DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668,  bigaddress340, Super_1_2_2_2);
WireDivision mux1_3_2_2(  DataOut31, DataOut33, DataOut35, DataOut37, DataOut39, DataOut41, DataOut43, DataOut45, DataOut47, DataOut49, DataOut51, DataOut53, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669,  bigaddress340, Super_1_3_2_2);
WireDivision mux1_4_2_2(  DataOut32, DataOut34, DataOut36, DataOut38, DataOut40, DataOut42, DataOut44, DataOut46, DataOut48, DataOut50, DataOut52, DataOut54, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut110, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670,  bigaddress340, Super_1_4_2_2);
WireDivision mux1_5_2_2(  DataOut33, DataOut35, DataOut37, DataOut39, DataOut41, DataOut43, DataOut45, DataOut47, DataOut49, DataOut51, DataOut53, DataOut55, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut111, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut167, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut223, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut279, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut335, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut391, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut447, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut503, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut559, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut615, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut671,  bigaddress340, Super_1_5_2_2);

WireDivision mux2_1_2_2(  DataOut57, DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut113, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut169, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut225, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut281, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut337, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut393, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut449, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut505, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut561, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut617, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut673, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695,  bigaddress340, Super_2_1_2_2);
WireDivision mux2_2_2_2(  DataOut58, DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696,  bigaddress340, Super_2_2_2_2);
WireDivision mux2_3_2_2(  DataOut59, DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut81, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697,  bigaddress340, Super_2_3_2_2);
WireDivision mux2_4_2_2(  DataOut60, DataOut62, DataOut64, DataOut66, DataOut68, DataOut70, DataOut72, DataOut74, DataOut76, DataOut78, DataOut80, DataOut82, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut138, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut194, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut250, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut306, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut362, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut418, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut474, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut530, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut586, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut642, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut698,  bigaddress340, Super_2_4_2_2);
WireDivision mux2_5_2_2(  DataOut61, DataOut63, DataOut65, DataOut67, DataOut69, DataOut71, DataOut73, DataOut75, DataOut77, DataOut79, DataOut81, DataOut83, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut139, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut195, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut251, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut307, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut363, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut419, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut475, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut531, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut587, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut643, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697, DataOut699,  bigaddress340, Super_2_5_2_2);

WireDivision mux3_1_2_2(  DataOut85, DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut141, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut197, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut253, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut309, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut365, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut421, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut477, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut533, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut589, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut645, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut701, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723,  bigaddress340, Super_3_1_2_2);
WireDivision mux3_2_2_2(  DataOut86, DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut702, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724,  bigaddress340, Super_3_2_2_2);
WireDivision mux3_3_2_2(  DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725,  bigaddress340, Super_3_3_2_2);
//WireDivision mux3_3_2_2(  DataOut87, DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725,  bigaddress340, Super_3_3_2_2);
WireDivision mux3_4_2_2(  DataOut88, DataOut90, DataOut92, DataOut94, DataOut96, DataOut98, DataOut100, DataOut102, DataOut104, DataOut106, DataOut108, DataOut110, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724, DataOut726,  bigaddress340, Super_3_4_2_2);
WireDivision mux3_5_2_2(  DataOut89, DataOut91, DataOut93, DataOut95, DataOut97, DataOut99, DataOut101, DataOut103, DataOut105, DataOut107, DataOut109, DataOut111, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut167, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut223, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut279, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut335, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut391, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut447, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut503, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut559, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut615, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut671, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725, DataOut727,  bigaddress340, Super_3_5_2_2);

WireDivision mux4_1_2_2(  DataOut113, DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut169, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut225, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut281, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut337, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut393, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut449, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut505, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut561, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut617, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut673, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut729, DataOut731, DataOut733, DataOut735, DataOut737, DataOut739, DataOut741, DataOut743, DataOut745, DataOut747, DataOut749, DataOut751,  bigaddress340, Super_4_1_2_2);
WireDivision mux4_2_2_2(  DataOut114, DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut170, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut226, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut282, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut338, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut394, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut450, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut506, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut562, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut618, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut674, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut730, DataOut732, DataOut734, DataOut736, DataOut738, DataOut740, DataOut742, DataOut744, DataOut746, DataOut748, DataOut750, DataOut752,  bigaddress340, Super_4_2_2_2);
WireDivision mux4_3_2_2(  DataOut115, DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut171, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut227, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut283, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut339, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut395, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut451, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut507, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut563, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut619, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut675, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697, DataOut731, DataOut733, DataOut735, DataOut737, DataOut739, DataOut741, DataOut743, DataOut745, DataOut747, DataOut749, DataOut751, DataOut753,  bigaddress340, Super_4_3_2_2);
WireDivision mux4_4_2_2(  DataOut116, DataOut118, DataOut120, DataOut122, DataOut124, DataOut126, DataOut128, DataOut130, DataOut132, DataOut134, DataOut136, DataOut138, DataOut172, DataOut174, DataOut176, DataOut178, DataOut180, DataOut182, DataOut184, DataOut186, DataOut188, DataOut190, DataOut192, DataOut194, DataOut228, DataOut230, DataOut232, DataOut234, DataOut236, DataOut238, DataOut240, DataOut242, DataOut244, DataOut246, DataOut248, DataOut250, DataOut284, DataOut286, DataOut288, DataOut290, DataOut292, DataOut294, DataOut296, DataOut298, DataOut300, DataOut302, DataOut304, DataOut306, DataOut340, DataOut342, DataOut344, DataOut346, DataOut348, DataOut350, DataOut352, DataOut354, DataOut356, DataOut358, DataOut360, DataOut362, DataOut396, DataOut398, DataOut400, DataOut402, DataOut404, DataOut406, DataOut408, DataOut410, DataOut412, DataOut414, DataOut416, DataOut418, DataOut452, DataOut454, DataOut456, DataOut458, DataOut460, DataOut462, DataOut464, DataOut466, DataOut468, DataOut470, DataOut472, DataOut474, DataOut508, DataOut510, DataOut512, DataOut514, DataOut516, DataOut518, DataOut520, DataOut522, DataOut524, DataOut526, DataOut528, DataOut530, DataOut564, DataOut566, DataOut568, DataOut570, DataOut572, DataOut574, DataOut576, DataOut578, DataOut580, DataOut582, DataOut584, DataOut586, DataOut620, DataOut622, DataOut624, DataOut626, DataOut628, DataOut630, DataOut632, DataOut634, DataOut636, DataOut638, DataOut640, DataOut642, DataOut676, DataOut678, DataOut680, DataOut682, DataOut684, DataOut686, DataOut688, DataOut690, DataOut692, DataOut694, DataOut696, DataOut698, DataOut732, DataOut734, DataOut736, DataOut738, DataOut740, DataOut742, DataOut744, DataOut746, DataOut748, DataOut750, DataOut752, DataOut754,  bigaddress340, Super_4_4_2_2);
WireDivision mux4_5_2_2(  DataOut117, DataOut119, DataOut121, DataOut123, DataOut125, DataOut127, DataOut129, DataOut131, DataOut133, DataOut135, DataOut137, DataOut139, DataOut173, DataOut175, DataOut177, DataOut179, DataOut181, DataOut183, DataOut185, DataOut187, DataOut189, DataOut191, DataOut193, DataOut195, DataOut229, DataOut231, DataOut233, DataOut235, DataOut237, DataOut239, DataOut241, DataOut243, DataOut245, DataOut247, DataOut249, DataOut251, DataOut285, DataOut287, DataOut289, DataOut291, DataOut293, DataOut295, DataOut297, DataOut299, DataOut301, DataOut303, DataOut305, DataOut307, DataOut341, DataOut343, DataOut345, DataOut347, DataOut349, DataOut351, DataOut353, DataOut355, DataOut357, DataOut359, DataOut361, DataOut363, DataOut397, DataOut399, DataOut401, DataOut403, DataOut405, DataOut407, DataOut409, DataOut411, DataOut413, DataOut415, DataOut417, DataOut419, DataOut453, DataOut455, DataOut457, DataOut459, DataOut461, DataOut463, DataOut465, DataOut467, DataOut469, DataOut471, DataOut473, DataOut475, DataOut509, DataOut511, DataOut513, DataOut515, DataOut517, DataOut519, DataOut521, DataOut523, DataOut525, DataOut527, DataOut529, DataOut531, DataOut565, DataOut567, DataOut569, DataOut571, DataOut573, DataOut575, DataOut577, DataOut579, DataOut581, DataOut583, DataOut585, DataOut587, DataOut621, DataOut623, DataOut625, DataOut627, DataOut629, DataOut631, DataOut633, DataOut635, DataOut637, DataOut639, DataOut641, DataOut643, DataOut677, DataOut679, DataOut681, DataOut683, DataOut685, DataOut687, DataOut689, DataOut691, DataOut693, DataOut695, DataOut697, DataOut699, DataOut733, DataOut735, DataOut737, DataOut739, DataOut741, DataOut743, DataOut745, DataOut747, DataOut749, DataOut751, DataOut753, DataOut755,  bigaddress340, Super_4_5_2_2);

WireDivision mux5_1_2_2(  DataOut141, DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut197, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut253, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut309, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut365, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut421, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut477, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut533, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut589, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut645, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut701, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut757, DataOut759, DataOut761, DataOut763, DataOut765, DataOut767, DataOut769, DataOut771, DataOut773, DataOut775, DataOut777, DataOut779,  bigaddress340, Super_5_1_2_2);
WireDivision mux5_2_2_2(  DataOut142, DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut198, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut254, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut310, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut366, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut422, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut478, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut534, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut590, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut646, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut702, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724, DataOut758, DataOut760, DataOut762, DataOut764, DataOut766, DataOut768, DataOut770, DataOut772, DataOut774, DataOut776, DataOut778, DataOut780,  bigaddress340, Super_5_2_2_2);
WireDivision mux5_3_2_2(  DataOut143, DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut199, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut255, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut311, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut367, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut423, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut479, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut535, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut591, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut647, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut703, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725, DataOut759, DataOut761, DataOut763, DataOut765, DataOut767, DataOut769, DataOut771, DataOut773, DataOut775, DataOut777, DataOut779, DataOut781,  bigaddress340, Super_5_3_2_2);
WireDivision mux5_4_2_2(  DataOut144, DataOut146, DataOut148, DataOut150, DataOut152, DataOut154, DataOut156, DataOut158, DataOut160, DataOut162, DataOut164, DataOut166, DataOut200, DataOut202, DataOut204, DataOut206, DataOut208, DataOut210, DataOut212, DataOut214, DataOut216, DataOut218, DataOut220, DataOut222, DataOut256, DataOut258, DataOut260, DataOut262, DataOut264, DataOut266, DataOut268, DataOut270, DataOut272, DataOut274, DataOut276, DataOut278, DataOut312, DataOut314, DataOut316, DataOut318, DataOut320, DataOut322, DataOut324, DataOut326, DataOut328, DataOut330, DataOut332, DataOut334, DataOut368, DataOut370, DataOut372, DataOut374, DataOut376, DataOut378, DataOut380, DataOut382, DataOut384, DataOut386, DataOut388, DataOut390, DataOut424, DataOut426, DataOut428, DataOut430, DataOut432, DataOut434, DataOut436, DataOut438, DataOut440, DataOut442, DataOut444, DataOut446, DataOut480, DataOut482, DataOut484, DataOut486, DataOut488, DataOut490, DataOut492, DataOut494, DataOut496, DataOut498, DataOut500, DataOut502, DataOut536, DataOut538, DataOut540, DataOut542, DataOut544, DataOut546, DataOut548, DataOut550, DataOut552, DataOut554, DataOut556, DataOut558, DataOut592, DataOut594, DataOut596, DataOut598, DataOut600, DataOut602, DataOut604, DataOut606, DataOut608, DataOut610, DataOut612, DataOut614, DataOut648, DataOut650, DataOut652, DataOut654, DataOut656, DataOut658, DataOut660, DataOut662, DataOut664, DataOut666, DataOut668, DataOut670, DataOut704, DataOut706, DataOut708, DataOut710, DataOut712, DataOut714, DataOut716, DataOut718, DataOut720, DataOut722, DataOut724, DataOut726, DataOut760, DataOut762, DataOut764, DataOut766, DataOut768, DataOut770, DataOut772, DataOut774, DataOut776, DataOut778, DataOut780, DataOut782,  bigaddress340, Super_5_4_2_2);
WireDivision mux5_5_2_2(  DataOut145, DataOut147, DataOut149, DataOut151, DataOut153, DataOut155, DataOut157, DataOut159, DataOut161, DataOut163, DataOut165, DataOut167, DataOut201, DataOut203, DataOut205, DataOut207, DataOut209, DataOut211, DataOut213, DataOut215, DataOut217, DataOut219, DataOut221, DataOut223, DataOut257, DataOut259, DataOut261, DataOut263, DataOut265, DataOut267, DataOut269, DataOut271, DataOut273, DataOut275, DataOut277, DataOut279, DataOut313, DataOut315, DataOut317, DataOut319, DataOut321, DataOut323, DataOut325, DataOut327, DataOut329, DataOut331, DataOut333, DataOut335, DataOut369, DataOut371, DataOut373, DataOut375, DataOut377, DataOut379, DataOut381, DataOut383, DataOut385, DataOut387, DataOut389, DataOut391, DataOut425, DataOut427, DataOut429, DataOut431, DataOut433, DataOut435, DataOut437, DataOut439, DataOut441, DataOut443, DataOut445, DataOut447, DataOut481, DataOut483, DataOut485, DataOut487, DataOut489, DataOut491, DataOut493, DataOut495, DataOut497, DataOut499, DataOut501, DataOut503, DataOut537, DataOut539, DataOut541, DataOut543, DataOut545, DataOut547, DataOut549, DataOut551, DataOut553, DataOut555, DataOut557, DataOut559, DataOut593, DataOut595, DataOut597, DataOut599, DataOut601, DataOut603, DataOut605, DataOut607, DataOut609, DataOut611, DataOut613, DataOut615, DataOut649, DataOut651, DataOut653, DataOut655, DataOut657, DataOut659, DataOut661, DataOut663, DataOut665, DataOut667, DataOut669, DataOut671, DataOut705, DataOut707, DataOut709, DataOut711, DataOut713, DataOut715, DataOut717, DataOut719, DataOut721, DataOut723, DataOut725, DataOut727, DataOut761, DataOut763, DataOut765, DataOut767, DataOut769, DataOut771, DataOut773, DataOut775, DataOut777, DataOut779, DataOut781, DataOut783,  bigaddress340, Super_5_5_2_2);



//----------------------------------------------------------------------------------------


MUX26X1_conv1 MUX1_1 ( Super_1_1_1_1 , Super_1_2_1_1 , Super_1_3_1_1 , Super_1_4_1_1 , Super_1_5_1_1 , Super_2_1_1_1 , Super_2_2_1_1 , Super_2_3_1_1 , Super_2_4_1_1 , Super_2_5_1_1 , Super_3_1_1_1 , Super_3_2_1_1 , Super_3_3_1_1 , Super_3_4_1_1 , Super_3_5_1_1 , Super_4_1_1_1 , Super_4_2_1_1 , Super_4_3_1_1 , Super_4_4_1_1 , Super_4_5_1_1 , Super_5_1_1_1 , Super_5_2_1_1 , Super_5_3_1_1 , Super_5_4_1_1 , Super_5_5_1_1 ,  DataOut784 , address , MUXout1_1 ); 
MUX26X1_conv1 MUX1_2 ( Super_1_1_1_2 , Super_1_2_1_2 , Super_1_3_1_2 , Super_1_4_1_2 , Super_1_5_1_2 , Super_2_1_1_2 , Super_2_2_1_2 , Super_2_3_1_2 , Super_2_4_1_2 , Super_2_5_1_2 , Super_3_1_1_2 , Super_3_2_1_2 , Super_3_3_1_2 , Super_3_4_1_2 , Super_3_5_1_2 , Super_4_1_1_2 , Super_4_2_1_2 , Super_4_3_1_2 , Super_4_4_1_2 , Super_4_5_1_2 , Super_5_1_1_2 , Super_5_2_1_2 , Super_5_3_1_2 , Super_5_4_1_2 , Super_5_5_1_2 ,  DataOut784 , address , MUXout1_2 ); 
MUX26X1_conv1 MUX2_1 ( Super_1_1_2_1 , Super_1_2_2_1 , Super_1_3_2_1 , Super_1_4_2_1 , Super_1_5_2_1 , Super_2_1_2_1 , Super_2_2_2_1 , Super_2_3_2_1 , Super_2_4_2_1 , Super_2_5_2_1 , Super_3_1_2_1 , Super_3_2_2_1 , Super_3_3_2_1 , Super_3_4_2_1 , Super_3_5_2_1 , Super_4_1_2_1 , Super_4_2_2_1 , Super_4_3_2_1 , Super_4_4_2_1 , Super_4_5_2_1 , Super_5_1_2_1 , Super_5_2_2_1 , Super_5_3_2_1 , Super_5_4_2_1 , Super_5_5_2_1 ,  DataOut784 , address , MUXout2_1 ); 
MUX26X1_conv1 MUX2_2 ( Super_1_1_2_2 , Super_1_2_2_2 , Super_1_3_2_2 , Super_1_4_2_2 , Super_1_5_2_2 , Super_2_1_2_2 , Super_2_2_2_2 , Super_2_3_2_2 , Super_2_4_2_2 , Super_2_5_2_2 , Super_3_1_2_2 , Super_3_2_2_2 , Super_3_3_2_2 , Super_3_4_2_2 , Super_3_5_2_2 , Super_4_1_2_2 , Super_4_2_2_2 , Super_4_3_2_2 , Super_4_4_2_2 , Super_4_5_2_2 , Super_5_1_2_2 , Super_5_2_2_2 , Super_5_3_2_2 , Super_5_4_2_2 , Super_5_5_2_2 ,  DataOut784 , address , MUXout2_2 ); 



MAC_26 MAC_F1_1_1  (ROMout1 , MUXout1_1  , clk , MACout_F1_1_1  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F1_1_2  (ROMout1 , MUXout1_2  , clk , MACout_F1_1_2  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F1_2_1  (ROMout1 , MUXout2_1  , clk , MACout_F1_2_1  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F1_2_2  (ROMout1 , MUXout2_2  , clk , MACout_F1_2_2  ,MAC_start, MAC_end , resetTheCounter);

MAC_26 MAC_F2_1_1  (ROMout2 , MUXout1_1  , clk , MACout_F2_1_1  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F2_1_2  (ROMout2 , MUXout1_2  , clk , MACout_F2_1_2  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F2_2_1  (ROMout2 , MUXout2_1  , clk , MACout_F2_2_1  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F2_2_2  (ROMout2 , MUXout2_2  , clk , MACout_F2_2_2  ,MAC_start, MAC_end , resetTheCounter);

MAC_26 MAC_F3_1_1  (ROMout3 , MUXout1_1  , clk , MACout_F3_1_1  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F3_1_2  (ROMout3 , MUXout1_2  , clk , MACout_F3_1_2  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F3_2_1  (ROMout3 , MUXout2_1  , clk , MACout_F3_2_1  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F3_2_2  (ROMout3 , MUXout2_2  , clk , MACout_F3_2_2  ,MAC_start, MAC_end , resetTheCounter);

MAC_26 MAC_F4_1_1  (ROMout4 , MUXout1_1  , clk , MACout_F4_1_1  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F4_1_2  (ROMout4 , MUXout1_2  , clk , MACout_F4_1_2  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F4_2_1  (ROMout4 , MUXout2_1  , clk , MACout_F4_2_1  ,MAC_start, MAC_end , resetTheCounter);
MAC_26 MAC_F4_2_2  (ROMout4 , MUXout2_2  , clk , MACout_F4_2_2  ,MAC_start, MAC_end , resetTheCounter);


RELU RELUF_1_1_1  ( MACout_F1_1_1  , clk , RELUout_F1_1_1  );
RELU RELUF_1_1_2  ( MACout_F1_1_2  , clk , RELUout_F1_1_2  );
RELU RELUF_1_2_1  ( MACout_F1_2_1  , clk , RELUout_F1_2_1  );
RELU RELUF_1_2_2  ( MACout_F1_2_2  , clk , RELUout_F1_2_2  ); 

RELU RELUF_2_1_1  ( MACout_F2_1_1  , clk , RELUout_F2_1_1  );
RELU RELUF_2_1_2  ( MACout_F2_1_2  , clk , RELUout_F2_1_2  );
RELU RELUF_2_2_1  ( MACout_F2_2_1  , clk , RELUout_F2_2_1  );
RELU RELUF_2_2_2  ( MACout_F2_2_2  , clk , RELUout_F2_2_2  );

RELU RELUF_3_1_1  ( MACout_F3_1_1  , clk , RELUout_F3_1_1  );
RELU RELUF_3_1_2  ( MACout_F3_1_2  , clk , RELUout_F3_1_2  );
RELU RELUF_3_2_1  ( MACout_F3_2_1  , clk , RELUout_F3_2_1  );
RELU RELUF_3_2_2  ( MACout_F3_2_2  , clk , RELUout_F3_2_2  );


RELU RELUF_4_1_1  ( MACout_F4_1_1  , clk , RELUout_F4_1_1  );
RELU RELUF_4_1_2  ( MACout_F4_1_2  , clk , RELUout_F4_1_2  );
RELU RELUF_4_2_1  ( MACout_F4_2_1  , clk , RELUout_F4_2_1  );
RELU RELUF_4_2_2  ( MACout_F4_2_2  , clk , RELUout_F4_2_2  );




/////

/*
OneRegister RAM_OUT_1_F1_1_1   ( clk , write2_1  , RELUout_F1_1_1  , Final_1_F1_1_1  );
OneRegister RAM_OUT_1_F1_1_2   ( clk , write2_1  , RELUout_F1_1_2  , Final_1_F1_1_2  );
OneRegister RAM_OUT_1_F1_2_1   ( clk , write2_1  , RELUout_F1_2_1  , Final_1_F1_2_1  );
OneRegister RAM_OUT_1_F1_2_2   ( clk , write2_1  , RELUout_F1_2_2  , Final_1_F1_2_2  );
OneRegister RAM_OUT_1_F2_1_1   ( clk , write2_1  , RELUout_F2_1_1  , Final_1_F2_1_1  );
OneRegister RAM_OUT_1_F2_1_2   ( clk , write2_1  , RELUout_F2_1_2  , Final_1_F2_1_2  );
OneRegister RAM_OUT_1_F2_2_1   ( clk , write2_1  , RELUout_F2_2_1  , Final_1_F2_2_1  );
OneRegister RAM_OUT_1_F2_2_2   ( clk , write2_1  , RELUout_F2_2_2  , Final_1_F2_2_2  );
OneRegister RAM_OUT_1_F3_1_1   ( clk , write2_1  , RELUout_F3_1_1  , Final_1_F3_1_1  );
OneRegister RAM_OUT_1_F3_1_2   ( clk , write2_1  , RELUout_F3_1_2  , Final_1_F3_1_2  );
OneRegister RAM_OUT_1_F3_2_1   ( clk , write2_1  , RELUout_F3_2_1  , Final_1_F3_2_1  );
OneRegister RAM_OUT_1_F3_2_2   ( clk , write2_1  , RELUout_F3_2_2  , Final_1_F3_2_2  );
OneRegister RAM_OUT_1_F4_1_1   ( clk , write2_1  , RELUout_F4_1_1  , Final_1_F4_1_1  );
OneRegister RAM_OUT_1_F4_1_2   ( clk , write2_1  , RELUout_F4_1_2  , Final_1_F4_1_2  );
OneRegister RAM_OUT_1_F4_2_1   ( clk , write2_1  , RELUout_F4_2_1  , Final_1_F4_2_1  );
OneRegister RAM_OUT_1_F4_2_2   ( clk , write2_1  , RELUout_F4_2_2  , Final_1_F4_2_2  );
OneRegister RAM_OUT_2_F1_1_1   ( clk , write2_2  , RELUout_F1_1_1  , Final_2_F1_1_1  );
OneRegister RAM_OUT_2_F1_1_2   ( clk , write2_2  , RELUout_F1_1_2  , Final_2_F1_1_2  );
OneRegister RAM_OUT_2_F1_2_1   ( clk , write2_2  , RELUout_F1_2_1  , Final_2_F1_2_1  );
OneRegister RAM_OUT_2_F1_2_2   ( clk , write2_2  , RELUout_F1_2_2  , Final_2_F1_2_2  );
OneRegister RAM_OUT_2_F2_1_1   ( clk , write2_2  , RELUout_F2_1_1  , Final_2_F2_1_1  );
OneRegister RAM_OUT_2_F2_1_2   ( clk , write2_2  , RELUout_F2_1_2  , Final_2_F2_1_2  );
OneRegister RAM_OUT_2_F2_2_1   ( clk , write2_2  , RELUout_F2_2_1  , Final_2_F2_2_1  );
OneRegister RAM_OUT_2_F2_2_2   ( clk , write2_2  , RELUout_F2_2_2  , Final_2_F2_2_2  );
OneRegister RAM_OUT_2_F3_1_1   ( clk , write2_2  , RELUout_F3_1_1  , Final_2_F3_1_1  );
OneRegister RAM_OUT_2_F3_1_2   ( clk , write2_2  , RELUout_F3_1_2  , Final_2_F3_1_2  );
OneRegister RAM_OUT_2_F3_2_1   ( clk , write2_2  , RELUout_F3_2_1  , Final_2_F3_2_1  );
OneRegister RAM_OUT_2_F3_2_2   ( clk , write2_2  , RELUout_F3_2_2  , Final_2_F3_2_2  );
OneRegister RAM_OUT_2_F4_1_1   ( clk , write2_2  , RELUout_F4_1_1  , Final_2_F4_1_1  );
OneRegister RAM_OUT_2_F4_1_2   ( clk , write2_2  , RELUout_F4_1_2  , Final_2_F4_1_2  );
OneRegister RAM_OUT_2_F4_2_1   ( clk , write2_2  , RELUout_F4_2_1  , Final_2_F4_2_1  );
OneRegister RAM_OUT_2_F4_2_2   ( clk , write2_2  , RELUout_F4_2_2  , Final_2_F4_2_2  );
OneRegister RAM_OUT_3_F1_1_1   ( clk , write2_3  , RELUout_F1_1_1  , Final_3_F1_1_1  );
OneRegister RAM_OUT_3_F1_1_2   ( clk , write2_3  , RELUout_F1_1_2  , Final_3_F1_1_2  );
OneRegister RAM_OUT_3_F1_2_1   ( clk , write2_3  , RELUout_F1_2_1  , Final_3_F1_2_1  );
OneRegister RAM_OUT_3_F1_2_2   ( clk , write2_3  , RELUout_F1_2_2  , Final_3_F1_2_2  );
OneRegister RAM_OUT_3_F2_1_1   ( clk , write2_3  , RELUout_F2_1_1  , Final_3_F2_1_1  );
OneRegister RAM_OUT_3_F2_1_2   ( clk , write2_3  , RELUout_F2_1_2  , Final_3_F2_1_2  );
OneRegister RAM_OUT_3_F2_2_1   ( clk , write2_3  , RELUout_F2_2_1  , Final_3_F2_2_1  );
OneRegister RAM_OUT_3_F2_2_2   ( clk , write2_3  , RELUout_F2_2_2  , Final_3_F2_2_2  );
OneRegister RAM_OUT_3_F3_1_1   ( clk , write2_3  , RELUout_F3_1_1  , Final_3_F3_1_1  );
OneRegister RAM_OUT_3_F3_1_2   ( clk , write2_3  , RELUout_F3_1_2  , Final_3_F3_1_2  );
OneRegister RAM_OUT_3_F3_2_1   ( clk , write2_3  , RELUout_F3_2_1  , Final_3_F3_2_1  );
OneRegister RAM_OUT_3_F3_2_2   ( clk , write2_3  , RELUout_F3_2_2  , Final_3_F3_2_2  );
OneRegister RAM_OUT_3_F4_1_1   ( clk , write2_3  , RELUout_F4_1_1  , Final_3_F4_1_1  );
OneRegister RAM_OUT_3_F4_1_2   ( clk , write2_3  , RELUout_F4_1_2  , Final_3_F4_1_2  );
OneRegister RAM_OUT_3_F4_2_1   ( clk , write2_3  , RELUout_F4_2_1  , Final_3_F4_2_1  );
OneRegister RAM_OUT_3_F4_2_2   ( clk , write2_3  , RELUout_F4_2_2  , Final_3_F4_2_2  );
OneRegister RAM_OUT_4_F1_1_1   ( clk , write2_4  , RELUout_F1_1_1  , Final_4_F1_1_1  );
OneRegister RAM_OUT_4_F1_1_2   ( clk , write2_4  , RELUout_F1_1_2  , Final_4_F1_1_2  );
OneRegister RAM_OUT_4_F1_2_1   ( clk , write2_4  , RELUout_F1_2_1  , Final_4_F1_2_1  );
OneRegister RAM_OUT_4_F1_2_2   ( clk , write2_4  , RELUout_F1_2_2  , Final_4_F1_2_2  );
OneRegister RAM_OUT_4_F2_1_1   ( clk , write2_4  , RELUout_F2_1_1  , Final_4_F2_1_1  );
OneRegister RAM_OUT_4_F2_1_2   ( clk , write2_4  , RELUout_F2_1_2  , Final_4_F2_1_2  );
OneRegister RAM_OUT_4_F2_2_1   ( clk , write2_4  , RELUout_F2_2_1  , Final_4_F2_2_1  );
OneRegister RAM_OUT_4_F2_2_2   ( clk , write2_4  , RELUout_F2_2_2  , Final_4_F2_2_2  );
OneRegister RAM_OUT_4_F3_1_1   ( clk , write2_4  , RELUout_F3_1_1  , Final_4_F3_1_1  );
OneRegister RAM_OUT_4_F3_1_2   ( clk , write2_4  , RELUout_F3_1_2  , Final_4_F3_1_2  );
OneRegister RAM_OUT_4_F3_2_1   ( clk , write2_4  , RELUout_F3_2_1  , Final_4_F3_2_1  );
OneRegister RAM_OUT_4_F3_2_2   ( clk , write2_4  , RELUout_F3_2_2  , Final_4_F3_2_2  );
OneRegister RAM_OUT_4_F4_1_1   ( clk , write2_4  , RELUout_F4_1_1  , Final_4_F4_1_1  );
OneRegister RAM_OUT_4_F4_1_2   ( clk , write2_4  , RELUout_F4_1_2  , Final_4_F4_1_2  );
OneRegister RAM_OUT_4_F4_2_1   ( clk , write2_4  , RELUout_F4_2_1  , Final_4_F4_2_1  );
OneRegister RAM_OUT_4_F4_2_2   ( clk , write2_4  , RELUout_F4_2_2  , Final_4_F4_2_2  );
OneRegister RAM_OUT_5_F1_1_1   ( clk , write2_5  , RELUout_F1_1_1  , Final_5_F1_1_1  );
OneRegister RAM_OUT_5_F1_1_2   ( clk , write2_5  , RELUout_F1_1_2  , Final_5_F1_1_2  );
OneRegister RAM_OUT_5_F1_2_1   ( clk , write2_5  , RELUout_F1_2_1  , Final_5_F1_2_1  );
OneRegister RAM_OUT_5_F1_2_2   ( clk , write2_5  , RELUout_F1_2_2  , Final_5_F1_2_2  );
OneRegister RAM_OUT_5_F2_1_1   ( clk , write2_5  , RELUout_F2_1_1  , Final_5_F2_1_1  );
OneRegister RAM_OUT_5_F2_1_2   ( clk , write2_5  , RELUout_F2_1_2  , Final_5_F2_1_2  );
OneRegister RAM_OUT_5_F2_2_1   ( clk , write2_5  , RELUout_F2_2_1  , Final_5_F2_2_1  );
OneRegister RAM_OUT_5_F2_2_2   ( clk , write2_5  , RELUout_F2_2_2  , Final_5_F2_2_2  );
OneRegister RAM_OUT_5_F3_1_1   ( clk , write2_5  , RELUout_F3_1_1  , Final_5_F3_1_1  );
OneRegister RAM_OUT_5_F3_1_2   ( clk , write2_5  , RELUout_F3_1_2  , Final_5_F3_1_2  );
OneRegister RAM_OUT_5_F3_2_1   ( clk , write2_5  , RELUout_F3_2_1  , Final_5_F3_2_1  );
OneRegister RAM_OUT_5_F3_2_2   ( clk , write2_5  , RELUout_F3_2_2  , Final_5_F3_2_2  );
OneRegister RAM_OUT_5_F4_1_1   ( clk , write2_5  , RELUout_F4_1_1  , Final_5_F4_1_1  );
OneRegister RAM_OUT_5_F4_1_2   ( clk , write2_5  , RELUout_F4_1_2  , Final_5_F4_1_2  );
OneRegister RAM_OUT_5_F4_2_1   ( clk , write2_5  , RELUout_F4_2_1  , Final_5_F4_2_1  );
OneRegister RAM_OUT_5_F4_2_2   ( clk , write2_5  , RELUout_F4_2_2  , Final_5_F4_2_2  );
OneRegister RAM_OUT_6_F1_1_1   ( clk , write2_6  , RELUout_F1_1_1  , Final_6_F1_1_1  );
OneRegister RAM_OUT_6_F1_1_2   ( clk , write2_6  , RELUout_F1_1_2  , Final_6_F1_1_2  );
OneRegister RAM_OUT_6_F1_2_1   ( clk , write2_6  , RELUout_F1_2_1  , Final_6_F1_2_1  );
OneRegister RAM_OUT_6_F1_2_2   ( clk , write2_6  , RELUout_F1_2_2  , Final_6_F1_2_2  );
OneRegister RAM_OUT_6_F2_1_1   ( clk , write2_6  , RELUout_F2_1_1  , Final_6_F2_1_1  );
OneRegister RAM_OUT_6_F2_1_2   ( clk , write2_6  , RELUout_F2_1_2  , Final_6_F2_1_2  );
OneRegister RAM_OUT_6_F2_2_1   ( clk , write2_6  , RELUout_F2_2_1  , Final_6_F2_2_1  );
OneRegister RAM_OUT_6_F2_2_2   ( clk , write2_6  , RELUout_F2_2_2  , Final_6_F2_2_2  );
OneRegister RAM_OUT_6_F3_1_1   ( clk , write2_6  , RELUout_F3_1_1  , Final_6_F3_1_1  );
OneRegister RAM_OUT_6_F3_1_2   ( clk , write2_6  , RELUout_F3_1_2  , Final_6_F3_1_2  );
OneRegister RAM_OUT_6_F3_2_1   ( clk , write2_6  , RELUout_F3_2_1  , Final_6_F3_2_1  );
OneRegister RAM_OUT_6_F3_2_2   ( clk , write2_6  , RELUout_F3_2_2  , Final_6_F3_2_2  );
OneRegister RAM_OUT_6_F4_1_1   ( clk , write2_6  , RELUout_F4_1_1  , Final_6_F4_1_1  );
OneRegister RAM_OUT_6_F4_1_2   ( clk , write2_6  , RELUout_F4_1_2  , Final_6_F4_1_2  );
OneRegister RAM_OUT_6_F4_2_1   ( clk , write2_6  , RELUout_F4_2_1  , Final_6_F4_2_1  );
OneRegister RAM_OUT_6_F4_2_2   ( clk , write2_6  , RELUout_F4_2_2  , Final_6_F4_2_2  );
OneRegister RAM_OUT_7_F1_1_1   ( clk , write2_7  , RELUout_F1_1_1  , Final_7_F1_1_1  );
OneRegister RAM_OUT_7_F1_1_2   ( clk , write2_7  , RELUout_F1_1_2  , Final_7_F1_1_2  );
OneRegister RAM_OUT_7_F1_2_1   ( clk , write2_7  , RELUout_F1_2_1  , Final_7_F1_2_1  );
OneRegister RAM_OUT_7_F1_2_2   ( clk , write2_7  , RELUout_F1_2_2  , Final_7_F1_2_2  );
OneRegister RAM_OUT_7_F2_1_1   ( clk , write2_7  , RELUout_F2_1_1  , Final_7_F2_1_1  );
OneRegister RAM_OUT_7_F2_1_2   ( clk , write2_7  , RELUout_F2_1_2  , Final_7_F2_1_2  );
OneRegister RAM_OUT_7_F2_2_1   ( clk , write2_7  , RELUout_F2_2_1  , Final_7_F2_2_1  );
OneRegister RAM_OUT_7_F2_2_2   ( clk , write2_7  , RELUout_F2_2_2  , Final_7_F2_2_2  );
OneRegister RAM_OUT_7_F3_1_1   ( clk , write2_7  , RELUout_F3_1_1  , Final_7_F3_1_1  );
OneRegister RAM_OUT_7_F3_1_2   ( clk , write2_7  , RELUout_F3_1_2  , Final_7_F3_1_2  );
OneRegister RAM_OUT_7_F3_2_1   ( clk , write2_7  , RELUout_F3_2_1  , Final_7_F3_2_1  );
OneRegister RAM_OUT_7_F3_2_2   ( clk , write2_7  , RELUout_F3_2_2  , Final_7_F3_2_2  );
OneRegister RAM_OUT_7_F4_1_1   ( clk , write2_7  , RELUout_F4_1_1  , Final_7_F4_1_1  );
OneRegister RAM_OUT_7_F4_1_2   ( clk , write2_7  , RELUout_F4_1_2  , Final_7_F4_1_2  );
OneRegister RAM_OUT_7_F4_2_1   ( clk , write2_7  , RELUout_F4_2_1  , Final_7_F4_2_1  );
OneRegister RAM_OUT_7_F4_2_2   ( clk , write2_7  , RELUout_F4_2_2  , Final_7_F4_2_2  );
OneRegister RAM_OUT_8_F1_1_1   ( clk , write2_8  , RELUout_F1_1_1  , Final_8_F1_1_1  );
OneRegister RAM_OUT_8_F1_1_2   ( clk , write2_8  , RELUout_F1_1_2  , Final_8_F1_1_2  );
OneRegister RAM_OUT_8_F1_2_1   ( clk , write2_8  , RELUout_F1_2_1  , Final_8_F1_2_1  );
OneRegister RAM_OUT_8_F1_2_2   ( clk , write2_8  , RELUout_F1_2_2  , Final_8_F1_2_2  );
OneRegister RAM_OUT_8_F2_1_1   ( clk , write2_8  , RELUout_F2_1_1  , Final_8_F2_1_1  );
OneRegister RAM_OUT_8_F2_1_2   ( clk , write2_8  , RELUout_F2_1_2  , Final_8_F2_1_2  );
OneRegister RAM_OUT_8_F2_2_1   ( clk , write2_8  , RELUout_F2_2_1  , Final_8_F2_2_1  );
OneRegister RAM_OUT_8_F2_2_2   ( clk , write2_8  , RELUout_F2_2_2  , Final_8_F2_2_2  );
OneRegister RAM_OUT_8_F3_1_1   ( clk , write2_8  , RELUout_F3_1_1  , Final_8_F3_1_1  );
OneRegister RAM_OUT_8_F3_1_2   ( clk , write2_8  , RELUout_F3_1_2  , Final_8_F3_1_2  );
OneRegister RAM_OUT_8_F3_2_1   ( clk , write2_8  , RELUout_F3_2_1  , Final_8_F3_2_1  );
OneRegister RAM_OUT_8_F3_2_2   ( clk , write2_8  , RELUout_F3_2_2  , Final_8_F3_2_2  );
OneRegister RAM_OUT_8_F4_1_1   ( clk , write2_8  , RELUout_F4_1_1  , Final_8_F4_1_1  );
OneRegister RAM_OUT_8_F4_1_2   ( clk , write2_8  , RELUout_F4_1_2  , Final_8_F4_1_2  );
OneRegister RAM_OUT_8_F4_2_1   ( clk , write2_8  , RELUout_F4_2_1  , Final_8_F4_2_1  );
OneRegister RAM_OUT_8_F4_2_2   ( clk , write2_8  , RELUout_F4_2_2  , Final_8_F4_2_2  );
OneRegister RAM_OUT_9_F1_1_1   ( clk , write2_9  , RELUout_F1_1_1  , Final_9_F1_1_1  );
OneRegister RAM_OUT_9_F1_1_2   ( clk , write2_9  , RELUout_F1_1_2  , Final_9_F1_1_2  );
OneRegister RAM_OUT_9_F1_2_1   ( clk , write2_9  , RELUout_F1_2_1  , Final_9_F1_2_1  );
OneRegister RAM_OUT_9_F1_2_2   ( clk , write2_9  , RELUout_F1_2_2  , Final_9_F1_2_2  );
OneRegister RAM_OUT_9_F2_1_1   ( clk , write2_9  , RELUout_F2_1_1  , Final_9_F2_1_1  );
OneRegister RAM_OUT_9_F2_1_2   ( clk , write2_9  , RELUout_F2_1_2  , Final_9_F2_1_2  );
OneRegister RAM_OUT_9_F2_2_1   ( clk , write2_9  , RELUout_F2_2_1  , Final_9_F2_2_1  );
OneRegister RAM_OUT_9_F2_2_2   ( clk , write2_9  , RELUout_F2_2_2  , Final_9_F2_2_2  );
OneRegister RAM_OUT_9_F3_1_1   ( clk , write2_9  , RELUout_F3_1_1  , Final_9_F3_1_1  );
OneRegister RAM_OUT_9_F3_1_2   ( clk , write2_9  , RELUout_F3_1_2  , Final_9_F3_1_2  );
OneRegister RAM_OUT_9_F3_2_1   ( clk , write2_9  , RELUout_F3_2_1  , Final_9_F3_2_1  );
OneRegister RAM_OUT_9_F3_2_2   ( clk , write2_9  , RELUout_F3_2_2  , Final_9_F3_2_2  );
OneRegister RAM_OUT_9_F4_1_1   ( clk , write2_9  , RELUout_F4_1_1  , Final_9_F4_1_1  );
OneRegister RAM_OUT_9_F4_1_2   ( clk , write2_9  , RELUout_F4_1_2  , Final_9_F4_1_2  );
OneRegister RAM_OUT_9_F4_2_1   ( clk , write2_9  , RELUout_F4_2_1  , Final_9_F4_2_1  );
OneRegister RAM_OUT_9_F4_2_2   ( clk , write2_9  , RELUout_F4_2_2  , Final_9_F4_2_2  );
OneRegister RAM_OUT_10_F1_1_1   ( clk , write2_10  , RELUout_F1_1_1  , Final_10_F1_1_1  );
OneRegister RAM_OUT_10_F1_1_2   ( clk , write2_10  , RELUout_F1_1_2  , Final_10_F1_1_2  );
OneRegister RAM_OUT_10_F1_2_1   ( clk , write2_10  , RELUout_F1_2_1  , Final_10_F1_2_1  );
OneRegister RAM_OUT_10_F1_2_2   ( clk , write2_10  , RELUout_F1_2_2  , Final_10_F1_2_2  );
OneRegister RAM_OUT_10_F2_1_1   ( clk , write2_10  , RELUout_F2_1_1  , Final_10_F2_1_1  );
OneRegister RAM_OUT_10_F2_1_2   ( clk , write2_10  , RELUout_F2_1_2  , Final_10_F2_1_2  );
OneRegister RAM_OUT_10_F2_2_1   ( clk , write2_10  , RELUout_F2_2_1  , Final_10_F2_2_1  );
OneRegister RAM_OUT_10_F2_2_2   ( clk , write2_10  , RELUout_F2_2_2  , Final_10_F2_2_2  );
OneRegister RAM_OUT_10_F3_1_1   ( clk , write2_10  , RELUout_F3_1_1  , Final_10_F3_1_1  );
OneRegister RAM_OUT_10_F3_1_2   ( clk , write2_10  , RELUout_F3_1_2  , Final_10_F3_1_2  );
OneRegister RAM_OUT_10_F3_2_1   ( clk , write2_10  , RELUout_F3_2_1  , Final_10_F3_2_1  );
OneRegister RAM_OUT_10_F3_2_2   ( clk , write2_10  , RELUout_F3_2_2  , Final_10_F3_2_2  );
OneRegister RAM_OUT_10_F4_1_1   ( clk , write2_10  , RELUout_F4_1_1  , Final_10_F4_1_1  );
OneRegister RAM_OUT_10_F4_1_2   ( clk , write2_10  , RELUout_F4_1_2  , Final_10_F4_1_2  );
OneRegister RAM_OUT_10_F4_2_1   ( clk , write2_10  , RELUout_F4_2_1  , Final_10_F4_2_1  );
OneRegister RAM_OUT_10_F4_2_2   ( clk , write2_10  , RELUout_F4_2_2  , Final_10_F4_2_2  );
OneRegister RAM_OUT_11_F1_1_1   ( clk , write2_11  , RELUout_F1_1_1  , Final_11_F1_1_1  );
OneRegister RAM_OUT_11_F1_1_2   ( clk , write2_11  , RELUout_F1_1_2  , Final_11_F1_1_2  );
OneRegister RAM_OUT_11_F1_2_1   ( clk , write2_11  , RELUout_F1_2_1  , Final_11_F1_2_1  );
OneRegister RAM_OUT_11_F1_2_2   ( clk , write2_11  , RELUout_F1_2_2  , Final_11_F1_2_2  );
OneRegister RAM_OUT_11_F2_1_1   ( clk , write2_11  , RELUout_F2_1_1  , Final_11_F2_1_1  );
OneRegister RAM_OUT_11_F2_1_2   ( clk , write2_11  , RELUout_F2_1_2  , Final_11_F2_1_2  );
OneRegister RAM_OUT_11_F2_2_1   ( clk , write2_11  , RELUout_F2_2_1  , Final_11_F2_2_1  );
OneRegister RAM_OUT_11_F2_2_2   ( clk , write2_11  , RELUout_F2_2_2  , Final_11_F2_2_2  );
OneRegister RAM_OUT_11_F3_1_1   ( clk , write2_11  , RELUout_F3_1_1  , Final_11_F3_1_1  );
OneRegister RAM_OUT_11_F3_1_2   ( clk , write2_11  , RELUout_F3_1_2  , Final_11_F3_1_2  );
OneRegister RAM_OUT_11_F3_2_1   ( clk , write2_11  , RELUout_F3_2_1  , Final_11_F3_2_1  );
OneRegister RAM_OUT_11_F3_2_2   ( clk , write2_11  , RELUout_F3_2_2  , Final_11_F3_2_2  );
OneRegister RAM_OUT_11_F4_1_1   ( clk , write2_11  , RELUout_F4_1_1  , Final_11_F4_1_1  );
OneRegister RAM_OUT_11_F4_1_2   ( clk , write2_11  , RELUout_F4_1_2  , Final_11_F4_1_2  );
OneRegister RAM_OUT_11_F4_2_1   ( clk , write2_11  , RELUout_F4_2_1  , Final_11_F4_2_1  );
OneRegister RAM_OUT_11_F4_2_2   ( clk , write2_11  , RELUout_F4_2_2  , Final_11_F4_2_2  );
OneRegister RAM_OUT_12_F1_1_1   ( clk , write2_12  , RELUout_F1_1_1  , Final_12_F1_1_1  );
OneRegister RAM_OUT_12_F1_1_2   ( clk , write2_12  , RELUout_F1_1_2  , Final_12_F1_1_2  );
OneRegister RAM_OUT_12_F1_2_1   ( clk , write2_12  , RELUout_F1_2_1  , Final_12_F1_2_1  );
OneRegister RAM_OUT_12_F1_2_2   ( clk , write2_12  , RELUout_F1_2_2  , Final_12_F1_2_2  );
OneRegister RAM_OUT_12_F2_1_1   ( clk , write2_12  , RELUout_F2_1_1  , Final_12_F2_1_1  );
OneRegister RAM_OUT_12_F2_1_2   ( clk , write2_12  , RELUout_F2_1_2  , Final_12_F2_1_2  );
OneRegister RAM_OUT_12_F2_2_1   ( clk , write2_12  , RELUout_F2_2_1  , Final_12_F2_2_1  );
OneRegister RAM_OUT_12_F2_2_2   ( clk , write2_12  , RELUout_F2_2_2  , Final_12_F2_2_2  );
OneRegister RAM_OUT_12_F3_1_1   ( clk , write2_12  , RELUout_F3_1_1  , Final_12_F3_1_1  );
OneRegister RAM_OUT_12_F3_1_2   ( clk , write2_12  , RELUout_F3_1_2  , Final_12_F3_1_2  );
OneRegister RAM_OUT_12_F3_2_1   ( clk , write2_12  , RELUout_F3_2_1  , Final_12_F3_2_1  );
OneRegister RAM_OUT_12_F3_2_2   ( clk , write2_12  , RELUout_F3_2_2  , Final_12_F3_2_2  );
OneRegister RAM_OUT_12_F4_1_1   ( clk , write2_12  , RELUout_F4_1_1  , Final_12_F4_1_1  );
OneRegister RAM_OUT_12_F4_1_2   ( clk , write2_12  , RELUout_F4_1_2  , Final_12_F4_1_2  );
OneRegister RAM_OUT_12_F4_2_1   ( clk , write2_12  , RELUout_F4_2_1  , Final_12_F4_2_1  );
OneRegister RAM_OUT_12_F4_2_2   ( clk , write2_12  , RELUout_F4_2_2  , Final_12_F4_2_2  );
OneRegister RAM_OUT_13_F1_1_1   ( clk , write2_13  , RELUout_F1_1_1  , Final_13_F1_1_1  );
OneRegister RAM_OUT_13_F1_1_2   ( clk , write2_13  , RELUout_F1_1_2  , Final_13_F1_1_2  );
OneRegister RAM_OUT_13_F1_2_1   ( clk , write2_13  , RELUout_F1_2_1  , Final_13_F1_2_1  );
OneRegister RAM_OUT_13_F1_2_2   ( clk , write2_13  , RELUout_F1_2_2  , Final_13_F1_2_2  );
OneRegister RAM_OUT_13_F2_1_1   ( clk , write2_13  , RELUout_F2_1_1  , Final_13_F2_1_1  );
OneRegister RAM_OUT_13_F2_1_2   ( clk , write2_13  , RELUout_F2_1_2  , Final_13_F2_1_2  );
OneRegister RAM_OUT_13_F2_2_1   ( clk , write2_13  , RELUout_F2_2_1  , Final_13_F2_2_1  );
OneRegister RAM_OUT_13_F2_2_2   ( clk , write2_13  , RELUout_F2_2_2  , Final_13_F2_2_2  );
OneRegister RAM_OUT_13_F3_1_1   ( clk , write2_13  , RELUout_F3_1_1  , Final_13_F3_1_1  );
OneRegister RAM_OUT_13_F3_1_2   ( clk , write2_13  , RELUout_F3_1_2  , Final_13_F3_1_2  );
OneRegister RAM_OUT_13_F3_2_1   ( clk , write2_13  , RELUout_F3_2_1  , Final_13_F3_2_1  );
OneRegister RAM_OUT_13_F3_2_2   ( clk , write2_13  , RELUout_F3_2_2  , Final_13_F3_2_2  );
OneRegister RAM_OUT_13_F4_1_1   ( clk , write2_13  , RELUout_F4_1_1  , Final_13_F4_1_1  );
OneRegister RAM_OUT_13_F4_1_2   ( clk , write2_13  , RELUout_F4_1_2  , Final_13_F4_1_2  );
OneRegister RAM_OUT_13_F4_2_1   ( clk , write2_13  , RELUout_F4_2_1  , Final_13_F4_2_1  );
OneRegister RAM_OUT_13_F4_2_2   ( clk , write2_13  , RELUout_F4_2_2  , Final_13_F4_2_2  );
OneRegister RAM_OUT_14_F1_1_1   ( clk , write2_14  , RELUout_F1_1_1  , Final_14_F1_1_1  );
OneRegister RAM_OUT_14_F1_1_2   ( clk , write2_14  , RELUout_F1_1_2  , Final_14_F1_1_2  );
OneRegister RAM_OUT_14_F1_2_1   ( clk , write2_14  , RELUout_F1_2_1  , Final_14_F1_2_1  );
OneRegister RAM_OUT_14_F1_2_2   ( clk , write2_14  , RELUout_F1_2_2  , Final_14_F1_2_2  );
OneRegister RAM_OUT_14_F2_1_1   ( clk , write2_14  , RELUout_F2_1_1  , Final_14_F2_1_1  );
OneRegister RAM_OUT_14_F2_1_2   ( clk , write2_14  , RELUout_F2_1_2  , Final_14_F2_1_2  );
OneRegister RAM_OUT_14_F2_2_1   ( clk , write2_14  , RELUout_F2_2_1  , Final_14_F2_2_1  );
OneRegister RAM_OUT_14_F2_2_2   ( clk , write2_14  , RELUout_F2_2_2  , Final_14_F2_2_2  );
OneRegister RAM_OUT_14_F3_1_1   ( clk , write2_14  , RELUout_F3_1_1  , Final_14_F3_1_1  );
OneRegister RAM_OUT_14_F3_1_2   ( clk , write2_14  , RELUout_F3_1_2  , Final_14_F3_1_2  );
OneRegister RAM_OUT_14_F3_2_1   ( clk , write2_14  , RELUout_F3_2_1  , Final_14_F3_2_1  );
OneRegister RAM_OUT_14_F3_2_2   ( clk , write2_14  , RELUout_F3_2_2  , Final_14_F3_2_2  );
OneRegister RAM_OUT_14_F4_1_1   ( clk , write2_14  , RELUout_F4_1_1  , Final_14_F4_1_1  );
OneRegister RAM_OUT_14_F4_1_2   ( clk , write2_14  , RELUout_F4_1_2  , Final_14_F4_1_2  );
OneRegister RAM_OUT_14_F4_2_1   ( clk , write2_14  , RELUout_F4_2_1  , Final_14_F4_2_1  );
OneRegister RAM_OUT_14_F4_2_2   ( clk , write2_14  , RELUout_F4_2_2  , Final_14_F4_2_2  );
OneRegister RAM_OUT_15_F1_1_1   ( clk , write2_15  , RELUout_F1_1_1  , Final_15_F1_1_1  );
OneRegister RAM_OUT_15_F1_1_2   ( clk , write2_15  , RELUout_F1_1_2  , Final_15_F1_1_2  );
OneRegister RAM_OUT_15_F1_2_1   ( clk , write2_15  , RELUout_F1_2_1  , Final_15_F1_2_1  );
OneRegister RAM_OUT_15_F1_2_2   ( clk , write2_15  , RELUout_F1_2_2  , Final_15_F1_2_2  );
OneRegister RAM_OUT_15_F2_1_1   ( clk , write2_15  , RELUout_F2_1_1  , Final_15_F2_1_1  );
OneRegister RAM_OUT_15_F2_1_2   ( clk , write2_15  , RELUout_F2_1_2  , Final_15_F2_1_2  );
OneRegister RAM_OUT_15_F2_2_1   ( clk , write2_15  , RELUout_F2_2_1  , Final_15_F2_2_1  );
OneRegister RAM_OUT_15_F2_2_2   ( clk , write2_15  , RELUout_F2_2_2  , Final_15_F2_2_2  );
OneRegister RAM_OUT_15_F3_1_1   ( clk , write2_15  , RELUout_F3_1_1  , Final_15_F3_1_1  );
OneRegister RAM_OUT_15_F3_1_2   ( clk , write2_15  , RELUout_F3_1_2  , Final_15_F3_1_2  );
OneRegister RAM_OUT_15_F3_2_1   ( clk , write2_15  , RELUout_F3_2_1  , Final_15_F3_2_1  );
OneRegister RAM_OUT_15_F3_2_2   ( clk , write2_15  , RELUout_F3_2_2  , Final_15_F3_2_2  );
OneRegister RAM_OUT_15_F4_1_1   ( clk , write2_15  , RELUout_F4_1_1  , Final_15_F4_1_1  );
OneRegister RAM_OUT_15_F4_1_2   ( clk , write2_15  , RELUout_F4_1_2  , Final_15_F4_1_2  );
OneRegister RAM_OUT_15_F4_2_1   ( clk , write2_15  , RELUout_F4_2_1  , Final_15_F4_2_1  );
OneRegister RAM_OUT_15_F4_2_2   ( clk , write2_15  , RELUout_F4_2_2  , Final_15_F4_2_2  );
OneRegister RAM_OUT_16_F1_1_1   ( clk , write2_16  , RELUout_F1_1_1  , Final_16_F1_1_1  );
OneRegister RAM_OUT_16_F1_1_2   ( clk , write2_16  , RELUout_F1_1_2  , Final_16_F1_1_2  );
OneRegister RAM_OUT_16_F1_2_1   ( clk , write2_16  , RELUout_F1_2_1  , Final_16_F1_2_1  );
OneRegister RAM_OUT_16_F1_2_2   ( clk , write2_16  , RELUout_F1_2_2  , Final_16_F1_2_2  );
OneRegister RAM_OUT_16_F2_1_1   ( clk , write2_16  , RELUout_F2_1_1  , Final_16_F2_1_1  );
OneRegister RAM_OUT_16_F2_1_2   ( clk , write2_16  , RELUout_F2_1_2  , Final_16_F2_1_2  );
OneRegister RAM_OUT_16_F2_2_1   ( clk , write2_16  , RELUout_F2_2_1  , Final_16_F2_2_1  );
OneRegister RAM_OUT_16_F2_2_2   ( clk , write2_16  , RELUout_F2_2_2  , Final_16_F2_2_2  );
OneRegister RAM_OUT_16_F3_1_1   ( clk , write2_16  , RELUout_F3_1_1  , Final_16_F3_1_1  );
OneRegister RAM_OUT_16_F3_1_2   ( clk , write2_16  , RELUout_F3_1_2  , Final_16_F3_1_2  );
OneRegister RAM_OUT_16_F3_2_1   ( clk , write2_16  , RELUout_F3_2_1  , Final_16_F3_2_1  );
OneRegister RAM_OUT_16_F3_2_2   ( clk , write2_16  , RELUout_F3_2_2  , Final_16_F3_2_2  );
OneRegister RAM_OUT_16_F4_1_1   ( clk , write2_16  , RELUout_F4_1_1  , Final_16_F4_1_1  );
OneRegister RAM_OUT_16_F4_1_2   ( clk , write2_16  , RELUout_F4_1_2  , Final_16_F4_1_2  );
OneRegister RAM_OUT_16_F4_2_1   ( clk , write2_16  , RELUout_F4_2_1  , Final_16_F4_2_1  );
OneRegister RAM_OUT_16_F4_2_2   ( clk , write2_16  , RELUout_F4_2_2  , Final_16_F4_2_2  );
OneRegister RAM_OUT_17_F1_1_1   ( clk , write2_17  , RELUout_F1_1_1  , Final_17_F1_1_1  );
OneRegister RAM_OUT_17_F1_1_2   ( clk , write2_17  , RELUout_F1_1_2  , Final_17_F1_1_2  );
OneRegister RAM_OUT_17_F1_2_1   ( clk , write2_17  , RELUout_F1_2_1  , Final_17_F1_2_1  );
OneRegister RAM_OUT_17_F1_2_2   ( clk , write2_17  , RELUout_F1_2_2  , Final_17_F1_2_2  );
OneRegister RAM_OUT_17_F2_1_1   ( clk , write2_17  , RELUout_F2_1_1  , Final_17_F2_1_1  );
OneRegister RAM_OUT_17_F2_1_2   ( clk , write2_17  , RELUout_F2_1_2  , Final_17_F2_1_2  );
OneRegister RAM_OUT_17_F2_2_1   ( clk , write2_17  , RELUout_F2_2_1  , Final_17_F2_2_1  );
OneRegister RAM_OUT_17_F2_2_2   ( clk , write2_17  , RELUout_F2_2_2  , Final_17_F2_2_2  );
OneRegister RAM_OUT_17_F3_1_1   ( clk , write2_17  , RELUout_F3_1_1  , Final_17_F3_1_1  );
OneRegister RAM_OUT_17_F3_1_2   ( clk , write2_17  , RELUout_F3_1_2  , Final_17_F3_1_2  );
OneRegister RAM_OUT_17_F3_2_1   ( clk , write2_17  , RELUout_F3_2_1  , Final_17_F3_2_1  );
OneRegister RAM_OUT_17_F3_2_2   ( clk , write2_17  , RELUout_F3_2_2  , Final_17_F3_2_2  );
OneRegister RAM_OUT_17_F4_1_1   ( clk , write2_17  , RELUout_F4_1_1  , Final_17_F4_1_1  );
OneRegister RAM_OUT_17_F4_1_2   ( clk , write2_17  , RELUout_F4_1_2  , Final_17_F4_1_2  );
OneRegister RAM_OUT_17_F4_2_1   ( clk , write2_17  , RELUout_F4_2_1  , Final_17_F4_2_1  );
OneRegister RAM_OUT_17_F4_2_2   ( clk , write2_17  , RELUout_F4_2_2  , Final_17_F4_2_2  );
OneRegister RAM_OUT_18_F1_1_1   ( clk , write2_18  , RELUout_F1_1_1  , Final_18_F1_1_1  );
OneRegister RAM_OUT_18_F1_1_2   ( clk , write2_18  , RELUout_F1_1_2  , Final_18_F1_1_2  );
OneRegister RAM_OUT_18_F1_2_1   ( clk , write2_18  , RELUout_F1_2_1  , Final_18_F1_2_1  );
OneRegister RAM_OUT_18_F1_2_2   ( clk , write2_18  , RELUout_F1_2_2  , Final_18_F1_2_2  );
OneRegister RAM_OUT_18_F2_1_1   ( clk , write2_18  , RELUout_F2_1_1  , Final_18_F2_1_1  );
OneRegister RAM_OUT_18_F2_1_2   ( clk , write2_18  , RELUout_F2_1_2  , Final_18_F2_1_2  );
OneRegister RAM_OUT_18_F2_2_1   ( clk , write2_18  , RELUout_F2_2_1  , Final_18_F2_2_1  );
OneRegister RAM_OUT_18_F2_2_2   ( clk , write2_18  , RELUout_F2_2_2  , Final_18_F2_2_2  );
OneRegister RAM_OUT_18_F3_1_1   ( clk , write2_18  , RELUout_F3_1_1  , Final_18_F3_1_1  );
OneRegister RAM_OUT_18_F3_1_2   ( clk , write2_18  , RELUout_F3_1_2  , Final_18_F3_1_2  );
OneRegister RAM_OUT_18_F3_2_1   ( clk , write2_18  , RELUout_F3_2_1  , Final_18_F3_2_1  );
OneRegister RAM_OUT_18_F3_2_2   ( clk , write2_18  , RELUout_F3_2_2  , Final_18_F3_2_2  );
OneRegister RAM_OUT_18_F4_1_1   ( clk , write2_18  , RELUout_F4_1_1  , Final_18_F4_1_1  );
OneRegister RAM_OUT_18_F4_1_2   ( clk , write2_18  , RELUout_F4_1_2  , Final_18_F4_1_2  );
OneRegister RAM_OUT_18_F4_2_1   ( clk , write2_18  , RELUout_F4_2_1  , Final_18_F4_2_1  );
OneRegister RAM_OUT_18_F4_2_2   ( clk , write2_18  , RELUout_F4_2_2  , Final_18_F4_2_2  );
OneRegister RAM_OUT_19_F1_1_1   ( clk , write2_19  , RELUout_F1_1_1  , Final_19_F1_1_1  );
OneRegister RAM_OUT_19_F1_1_2   ( clk , write2_19  , RELUout_F1_1_2  , Final_19_F1_1_2  );
OneRegister RAM_OUT_19_F1_2_1   ( clk , write2_19  , RELUout_F1_2_1  , Final_19_F1_2_1  );
OneRegister RAM_OUT_19_F1_2_2   ( clk , write2_19  , RELUout_F1_2_2  , Final_19_F1_2_2  );
OneRegister RAM_OUT_19_F2_1_1   ( clk , write2_19  , RELUout_F2_1_1  , Final_19_F2_1_1  );
OneRegister RAM_OUT_19_F2_1_2   ( clk , write2_19  , RELUout_F2_1_2  , Final_19_F2_1_2  );
OneRegister RAM_OUT_19_F2_2_1   ( clk , write2_19  , RELUout_F2_2_1  , Final_19_F2_2_1  );
OneRegister RAM_OUT_19_F2_2_2   ( clk , write2_19  , RELUout_F2_2_2  , Final_19_F2_2_2  );
OneRegister RAM_OUT_19_F3_1_1   ( clk , write2_19  , RELUout_F3_1_1  , Final_19_F3_1_1  );
OneRegister RAM_OUT_19_F3_1_2   ( clk , write2_19  , RELUout_F3_1_2  , Final_19_F3_1_2  );
OneRegister RAM_OUT_19_F3_2_1   ( clk , write2_19  , RELUout_F3_2_1  , Final_19_F3_2_1  );
OneRegister RAM_OUT_19_F3_2_2   ( clk , write2_19  , RELUout_F3_2_2  , Final_19_F3_2_2  );
OneRegister RAM_OUT_19_F4_1_1   ( clk , write2_19  , RELUout_F4_1_1  , Final_19_F4_1_1  );
OneRegister RAM_OUT_19_F4_1_2   ( clk , write2_19  , RELUout_F4_1_2  , Final_19_F4_1_2  );
OneRegister RAM_OUT_19_F4_2_1   ( clk , write2_19  , RELUout_F4_2_1  , Final_19_F4_2_1  );
OneRegister RAM_OUT_19_F4_2_2   ( clk , write2_19  , RELUout_F4_2_2  , Final_19_F4_2_2  );
OneRegister RAM_OUT_20_F1_1_1   ( clk , write2_20  , RELUout_F1_1_1  , Final_20_F1_1_1  );
OneRegister RAM_OUT_20_F1_1_2   ( clk , write2_20  , RELUout_F1_1_2  , Final_20_F1_1_2  );
OneRegister RAM_OUT_20_F1_2_1   ( clk , write2_20  , RELUout_F1_2_1  , Final_20_F1_2_1  );
OneRegister RAM_OUT_20_F1_2_2   ( clk , write2_20  , RELUout_F1_2_2  , Final_20_F1_2_2  );
OneRegister RAM_OUT_20_F2_1_1   ( clk , write2_20  , RELUout_F2_1_1  , Final_20_F2_1_1  );
OneRegister RAM_OUT_20_F2_1_2   ( clk , write2_20  , RELUout_F2_1_2  , Final_20_F2_1_2  );
OneRegister RAM_OUT_20_F2_2_1   ( clk , write2_20  , RELUout_F2_2_1  , Final_20_F2_2_1  );
OneRegister RAM_OUT_20_F2_2_2   ( clk , write2_20  , RELUout_F2_2_2  , Final_20_F2_2_2  );
OneRegister RAM_OUT_20_F3_1_1   ( clk , write2_20  , RELUout_F3_1_1  , Final_20_F3_1_1  );
OneRegister RAM_OUT_20_F3_1_2   ( clk , write2_20  , RELUout_F3_1_2  , Final_20_F3_1_2  );
OneRegister RAM_OUT_20_F3_2_1   ( clk , write2_20  , RELUout_F3_2_1  , Final_20_F3_2_1  );
OneRegister RAM_OUT_20_F3_2_2   ( clk , write2_20  , RELUout_F3_2_2  , Final_20_F3_2_2  );
OneRegister RAM_OUT_20_F4_1_1   ( clk , write2_20  , RELUout_F4_1_1  , Final_20_F4_1_1  );
OneRegister RAM_OUT_20_F4_1_2   ( clk , write2_20  , RELUout_F4_1_2  , Final_20_F4_1_2  );
OneRegister RAM_OUT_20_F4_2_1   ( clk , write2_20  , RELUout_F4_2_1  , Final_20_F4_2_1  );
OneRegister RAM_OUT_20_F4_2_2   ( clk , write2_20  , RELUout_F4_2_2  , Final_20_F4_2_2  );
OneRegister RAM_OUT_21_F1_1_1   ( clk , write2_21  , RELUout_F1_1_1  , Final_21_F1_1_1  );
OneRegister RAM_OUT_21_F1_1_2   ( clk , write2_21  , RELUout_F1_1_2  , Final_21_F1_1_2  );
OneRegister RAM_OUT_21_F1_2_1   ( clk , write2_21  , RELUout_F1_2_1  , Final_21_F1_2_1  );
OneRegister RAM_OUT_21_F1_2_2   ( clk , write2_21  , RELUout_F1_2_2  , Final_21_F1_2_2  );
OneRegister RAM_OUT_21_F2_1_1   ( clk , write2_21  , RELUout_F2_1_1  , Final_21_F2_1_1  );
OneRegister RAM_OUT_21_F2_1_2   ( clk , write2_21  , RELUout_F2_1_2  , Final_21_F2_1_2  );
OneRegister RAM_OUT_21_F2_2_1   ( clk , write2_21  , RELUout_F2_2_1  , Final_21_F2_2_1  );
OneRegister RAM_OUT_21_F2_2_2   ( clk , write2_21  , RELUout_F2_2_2  , Final_21_F2_2_2  );
OneRegister RAM_OUT_21_F3_1_1   ( clk , write2_21  , RELUout_F3_1_1  , Final_21_F3_1_1  );
OneRegister RAM_OUT_21_F3_1_2   ( clk , write2_21  , RELUout_F3_1_2  , Final_21_F3_1_2  );
OneRegister RAM_OUT_21_F3_2_1   ( clk , write2_21  , RELUout_F3_2_1  , Final_21_F3_2_1  );
OneRegister RAM_OUT_21_F3_2_2   ( clk , write2_21  , RELUout_F3_2_2  , Final_21_F3_2_2  );
OneRegister RAM_OUT_21_F4_1_1   ( clk , write2_21  , RELUout_F4_1_1  , Final_21_F4_1_1  );
OneRegister RAM_OUT_21_F4_1_2   ( clk , write2_21  , RELUout_F4_1_2  , Final_21_F4_1_2  );
OneRegister RAM_OUT_21_F4_2_1   ( clk , write2_21  , RELUout_F4_2_1  , Final_21_F4_2_1  );
OneRegister RAM_OUT_21_F4_2_2   ( clk , write2_21  , RELUout_F4_2_2  , Final_21_F4_2_2  );
OneRegister RAM_OUT_22_F1_1_1   ( clk , write2_22  , RELUout_F1_1_1  , Final_22_F1_1_1  );
OneRegister RAM_OUT_22_F1_1_2   ( clk , write2_22  , RELUout_F1_1_2  , Final_22_F1_1_2  );
OneRegister RAM_OUT_22_F1_2_1   ( clk , write2_22  , RELUout_F1_2_1  , Final_22_F1_2_1  );
OneRegister RAM_OUT_22_F1_2_2   ( clk , write2_22  , RELUout_F1_2_2  , Final_22_F1_2_2  );
OneRegister RAM_OUT_22_F2_1_1   ( clk , write2_22  , RELUout_F2_1_1  , Final_22_F2_1_1  );
OneRegister RAM_OUT_22_F2_1_2   ( clk , write2_22  , RELUout_F2_1_2  , Final_22_F2_1_2  );
OneRegister RAM_OUT_22_F2_2_1   ( clk , write2_22  , RELUout_F2_2_1  , Final_22_F2_2_1  );
OneRegister RAM_OUT_22_F2_2_2   ( clk , write2_22  , RELUout_F2_2_2  , Final_22_F2_2_2  );
OneRegister RAM_OUT_22_F3_1_1   ( clk , write2_22  , RELUout_F3_1_1  , Final_22_F3_1_1  );
OneRegister RAM_OUT_22_F3_1_2   ( clk , write2_22  , RELUout_F3_1_2  , Final_22_F3_1_2  );
OneRegister RAM_OUT_22_F3_2_1   ( clk , write2_22  , RELUout_F3_2_1  , Final_22_F3_2_1  );
OneRegister RAM_OUT_22_F3_2_2   ( clk , write2_22  , RELUout_F3_2_2  , Final_22_F3_2_2  );
OneRegister RAM_OUT_22_F4_1_1   ( clk , write2_22  , RELUout_F4_1_1  , Final_22_F4_1_1  );
OneRegister RAM_OUT_22_F4_1_2   ( clk , write2_22  , RELUout_F4_1_2  , Final_22_F4_1_2  );
OneRegister RAM_OUT_22_F4_2_1   ( clk , write2_22  , RELUout_F4_2_1  , Final_22_F4_2_1  );
OneRegister RAM_OUT_22_F4_2_2   ( clk , write2_22  , RELUout_F4_2_2  , Final_22_F4_2_2  );
OneRegister RAM_OUT_23_F1_1_1   ( clk , write2_23  , RELUout_F1_1_1  , Final_23_F1_1_1  );
OneRegister RAM_OUT_23_F1_1_2   ( clk , write2_23  , RELUout_F1_1_2  , Final_23_F1_1_2  );
OneRegister RAM_OUT_23_F1_2_1   ( clk , write2_23  , RELUout_F1_2_1  , Final_23_F1_2_1  );
OneRegister RAM_OUT_23_F1_2_2   ( clk , write2_23  , RELUout_F1_2_2  , Final_23_F1_2_2  );
OneRegister RAM_OUT_23_F2_1_1   ( clk , write2_23  , RELUout_F2_1_1  , Final_23_F2_1_1  );
OneRegister RAM_OUT_23_F2_1_2   ( clk , write2_23  , RELUout_F2_1_2  , Final_23_F2_1_2  );
OneRegister RAM_OUT_23_F2_2_1   ( clk , write2_23  , RELUout_F2_2_1  , Final_23_F2_2_1  );
OneRegister RAM_OUT_23_F2_2_2   ( clk , write2_23  , RELUout_F2_2_2  , Final_23_F2_2_2  );
OneRegister RAM_OUT_23_F3_1_1   ( clk , write2_23  , RELUout_F3_1_1  , Final_23_F3_1_1  );
OneRegister RAM_OUT_23_F3_1_2   ( clk , write2_23  , RELUout_F3_1_2  , Final_23_F3_1_2  );
OneRegister RAM_OUT_23_F3_2_1   ( clk , write2_23  , RELUout_F3_2_1  , Final_23_F3_2_1  );
OneRegister RAM_OUT_23_F3_2_2   ( clk , write2_23  , RELUout_F3_2_2  , Final_23_F3_2_2  );
OneRegister RAM_OUT_23_F4_1_1   ( clk , write2_23  , RELUout_F4_1_1  , Final_23_F4_1_1  );
OneRegister RAM_OUT_23_F4_1_2   ( clk , write2_23  , RELUout_F4_1_2  , Final_23_F4_1_2  );
OneRegister RAM_OUT_23_F4_2_1   ( clk , write2_23  , RELUout_F4_2_1  , Final_23_F4_2_1  );
OneRegister RAM_OUT_23_F4_2_2   ( clk , write2_23  , RELUout_F4_2_2  , Final_23_F4_2_2  );
OneRegister RAM_OUT_24_F1_1_1   ( clk , write2_24  , RELUout_F1_1_1  , Final_24_F1_1_1  );
OneRegister RAM_OUT_24_F1_1_2   ( clk , write2_24  , RELUout_F1_1_2  , Final_24_F1_1_2  );
OneRegister RAM_OUT_24_F1_2_1   ( clk , write2_24  , RELUout_F1_2_1  , Final_24_F1_2_1  );
OneRegister RAM_OUT_24_F1_2_2   ( clk , write2_24  , RELUout_F1_2_2  , Final_24_F1_2_2  );
OneRegister RAM_OUT_24_F2_1_1   ( clk , write2_24  , RELUout_F2_1_1  , Final_24_F2_1_1  );
OneRegister RAM_OUT_24_F2_1_2   ( clk , write2_24  , RELUout_F2_1_2  , Final_24_F2_1_2  );
OneRegister RAM_OUT_24_F2_2_1   ( clk , write2_24  , RELUout_F2_2_1  , Final_24_F2_2_1  );
OneRegister RAM_OUT_24_F2_2_2   ( clk , write2_24  , RELUout_F2_2_2  , Final_24_F2_2_2  );
OneRegister RAM_OUT_24_F3_1_1   ( clk , write2_24  , RELUout_F3_1_1  , Final_24_F3_1_1  );
OneRegister RAM_OUT_24_F3_1_2   ( clk , write2_24  , RELUout_F3_1_2  , Final_24_F3_1_2  );
OneRegister RAM_OUT_24_F3_2_1   ( clk , write2_24  , RELUout_F3_2_1  , Final_24_F3_2_1  );
OneRegister RAM_OUT_24_F3_2_2   ( clk , write2_24  , RELUout_F3_2_2  , Final_24_F3_2_2  );
OneRegister RAM_OUT_24_F4_1_1   ( clk , write2_24  , RELUout_F4_1_1  , Final_24_F4_1_1  );
OneRegister RAM_OUT_24_F4_1_2   ( clk , write2_24  , RELUout_F4_1_2  , Final_24_F4_1_2  );
OneRegister RAM_OUT_24_F4_2_1   ( clk , write2_24  , RELUout_F4_2_1  , Final_24_F4_2_1  );
OneRegister RAM_OUT_24_F4_2_2   ( clk , write2_24  , RELUout_F4_2_2  , Final_24_F4_2_2  );
OneRegister RAM_OUT_25_F1_1_1   ( clk , write2_25  , RELUout_F1_1_1  , Final_25_F1_1_1  );
OneRegister RAM_OUT_25_F1_1_2   ( clk , write2_25  , RELUout_F1_1_2  , Final_25_F1_1_2  );
OneRegister RAM_OUT_25_F1_2_1   ( clk , write2_25  , RELUout_F1_2_1  , Final_25_F1_2_1  );
OneRegister RAM_OUT_25_F1_2_2   ( clk , write2_25  , RELUout_F1_2_2  , Final_25_F1_2_2  );
OneRegister RAM_OUT_25_F2_1_1   ( clk , write2_25  , RELUout_F2_1_1  , Final_25_F2_1_1  );
OneRegister RAM_OUT_25_F2_1_2   ( clk , write2_25  , RELUout_F2_1_2  , Final_25_F2_1_2  );
OneRegister RAM_OUT_25_F2_2_1   ( clk , write2_25  , RELUout_F2_2_1  , Final_25_F2_2_1  );
OneRegister RAM_OUT_25_F2_2_2   ( clk , write2_25  , RELUout_F2_2_2  , Final_25_F2_2_2  );
OneRegister RAM_OUT_25_F3_1_1   ( clk , write2_25  , RELUout_F3_1_1  , Final_25_F3_1_1  );
OneRegister RAM_OUT_25_F3_1_2   ( clk , write2_25  , RELUout_F3_1_2  , Final_25_F3_1_2  );
OneRegister RAM_OUT_25_F3_2_1   ( clk , write2_25  , RELUout_F3_2_1  , Final_25_F3_2_1  );
OneRegister RAM_OUT_25_F3_2_2   ( clk , write2_25  , RELUout_F3_2_2  , Final_25_F3_2_2  );
OneRegister RAM_OUT_25_F4_1_1   ( clk , write2_25  , RELUout_F4_1_1  , Final_25_F4_1_1  );
OneRegister RAM_OUT_25_F4_1_2   ( clk , write2_25  , RELUout_F4_1_2  , Final_25_F4_1_2  );
OneRegister RAM_OUT_25_F4_2_1   ( clk , write2_25  , RELUout_F4_2_1  , Final_25_F4_2_1  );
OneRegister RAM_OUT_25_F4_2_2   ( clk , write2_25  , RELUout_F4_2_2  , Final_25_F4_2_2  );
OneRegister RAM_OUT_26_F1_1_1   ( clk , write2_26  , RELUout_F1_1_1  , Final_26_F1_1_1  );
OneRegister RAM_OUT_26_F1_1_2   ( clk , write2_26  , RELUout_F1_1_2  , Final_26_F1_1_2  );
OneRegister RAM_OUT_26_F1_2_1   ( clk , write2_26  , RELUout_F1_2_1  , Final_26_F1_2_1  );
OneRegister RAM_OUT_26_F1_2_2   ( clk , write2_26  , RELUout_F1_2_2  , Final_26_F1_2_2  );
OneRegister RAM_OUT_26_F2_1_1   ( clk , write2_26  , RELUout_F2_1_1  , Final_26_F2_1_1  );
OneRegister RAM_OUT_26_F2_1_2   ( clk , write2_26  , RELUout_F2_1_2  , Final_26_F2_1_2  );
OneRegister RAM_OUT_26_F2_2_1   ( clk , write2_26  , RELUout_F2_2_1  , Final_26_F2_2_1  );
OneRegister RAM_OUT_26_F2_2_2   ( clk , write2_26  , RELUout_F2_2_2  , Final_26_F2_2_2  );
OneRegister RAM_OUT_26_F3_1_1   ( clk , write2_26  , RELUout_F3_1_1  , Final_26_F3_1_1  );
OneRegister RAM_OUT_26_F3_1_2   ( clk , write2_26  , RELUout_F3_1_2  , Final_26_F3_1_2  );
OneRegister RAM_OUT_26_F3_2_1   ( clk , write2_26  , RELUout_F3_2_1  , Final_26_F3_2_1  );
OneRegister RAM_OUT_26_F3_2_2   ( clk , write2_26  , RELUout_F3_2_2  , Final_26_F3_2_2  );
OneRegister RAM_OUT_26_F4_1_1   ( clk , write2_26  , RELUout_F4_1_1  , Final_26_F4_1_1  );
OneRegister RAM_OUT_26_F4_1_2   ( clk , write2_26  , RELUout_F4_1_2  , Final_26_F4_1_2  );
OneRegister RAM_OUT_26_F4_2_1   ( clk , write2_26  , RELUout_F4_2_1  , Final_26_F4_2_1  );
OneRegister RAM_OUT_26_F4_2_2   ( clk , write2_26  , RELUout_F4_2_2  , Final_26_F4_2_2  );
OneRegister RAM_OUT_27_F1_1_1   ( clk , write2_27  , RELUout_F1_1_1  , Final_27_F1_1_1  );
OneRegister RAM_OUT_27_F1_1_2   ( clk , write2_27  , RELUout_F1_1_2  , Final_27_F1_1_2  );
OneRegister RAM_OUT_27_F1_2_1   ( clk , write2_27  , RELUout_F1_2_1  , Final_27_F1_2_1  );
OneRegister RAM_OUT_27_F1_2_2   ( clk , write2_27  , RELUout_F1_2_2  , Final_27_F1_2_2  );
OneRegister RAM_OUT_27_F2_1_1   ( clk , write2_27  , RELUout_F2_1_1  , Final_27_F2_1_1  );
OneRegister RAM_OUT_27_F2_1_2   ( clk , write2_27  , RELUout_F2_1_2  , Final_27_F2_1_2  );
OneRegister RAM_OUT_27_F2_2_1   ( clk , write2_27  , RELUout_F2_2_1  , Final_27_F2_2_1  );
OneRegister RAM_OUT_27_F2_2_2   ( clk , write2_27  , RELUout_F2_2_2  , Final_27_F2_2_2  );
OneRegister RAM_OUT_27_F3_1_1   ( clk , write2_27  , RELUout_F3_1_1  , Final_27_F3_1_1  );
OneRegister RAM_OUT_27_F3_1_2   ( clk , write2_27  , RELUout_F3_1_2  , Final_27_F3_1_2  );
OneRegister RAM_OUT_27_F3_2_1   ( clk , write2_27  , RELUout_F3_2_1  , Final_27_F3_2_1  );
OneRegister RAM_OUT_27_F3_2_2   ( clk , write2_27  , RELUout_F3_2_2  , Final_27_F3_2_2  );
OneRegister RAM_OUT_27_F4_1_1   ( clk , write2_27  , RELUout_F4_1_1  , Final_27_F4_1_1  );
OneRegister RAM_OUT_27_F4_1_2   ( clk , write2_27  , RELUout_F4_1_2  , Final_27_F4_1_2  );
OneRegister RAM_OUT_27_F4_2_1   ( clk , write2_27  , RELUout_F4_2_1  , Final_27_F4_2_1  );
OneRegister RAM_OUT_27_F4_2_2   ( clk , write2_27  , RELUout_F4_2_2  , Final_27_F4_2_2  );
OneRegister RAM_OUT_28_F1_1_1   ( clk , write2_28  , RELUout_F1_1_1  , Final_28_F1_1_1  );
OneRegister RAM_OUT_28_F1_1_2   ( clk , write2_28  , RELUout_F1_1_2  , Final_28_F1_1_2  );
OneRegister RAM_OUT_28_F1_2_1   ( clk , write2_28  , RELUout_F1_2_1  , Final_28_F1_2_1  );
OneRegister RAM_OUT_28_F1_2_2   ( clk , write2_28  , RELUout_F1_2_2  , Final_28_F1_2_2  );
OneRegister RAM_OUT_28_F2_1_1   ( clk , write2_28  , RELUout_F2_1_1  , Final_28_F2_1_1  );
OneRegister RAM_OUT_28_F2_1_2   ( clk , write2_28  , RELUout_F2_1_2  , Final_28_F2_1_2  );
OneRegister RAM_OUT_28_F2_2_1   ( clk , write2_28  , RELUout_F2_2_1  , Final_28_F2_2_1  );
OneRegister RAM_OUT_28_F2_2_2   ( clk , write2_28  , RELUout_F2_2_2  , Final_28_F2_2_2  );
OneRegister RAM_OUT_28_F3_1_1   ( clk , write2_28  , RELUout_F3_1_1  , Final_28_F3_1_1  );
OneRegister RAM_OUT_28_F3_1_2   ( clk , write2_28  , RELUout_F3_1_2  , Final_28_F3_1_2  );
OneRegister RAM_OUT_28_F3_2_1   ( clk , write2_28  , RELUout_F3_2_1  , Final_28_F3_2_1  );
OneRegister RAM_OUT_28_F3_2_2   ( clk , write2_28  , RELUout_F3_2_2  , Final_28_F3_2_2  );
OneRegister RAM_OUT_28_F4_1_1   ( clk , write2_28  , RELUout_F4_1_1  , Final_28_F4_1_1  );
OneRegister RAM_OUT_28_F4_1_2   ( clk , write2_28  , RELUout_F4_1_2  , Final_28_F4_1_2  );
OneRegister RAM_OUT_28_F4_2_1   ( clk , write2_28  , RELUout_F4_2_1  , Final_28_F4_2_1  );
OneRegister RAM_OUT_28_F4_2_2   ( clk , write2_28  , RELUout_F4_2_2  , Final_28_F4_2_2  );
OneRegister RAM_OUT_29_F1_1_1   ( clk , write2_29  , RELUout_F1_1_1  , Final_29_F1_1_1  );
OneRegister RAM_OUT_29_F1_1_2   ( clk , write2_29  , RELUout_F1_1_2  , Final_29_F1_1_2  );
OneRegister RAM_OUT_29_F1_2_1   ( clk , write2_29  , RELUout_F1_2_1  , Final_29_F1_2_1  );
OneRegister RAM_OUT_29_F1_2_2   ( clk , write2_29  , RELUout_F1_2_2  , Final_29_F1_2_2  );
OneRegister RAM_OUT_29_F2_1_1   ( clk , write2_29  , RELUout_F2_1_1  , Final_29_F2_1_1  );
OneRegister RAM_OUT_29_F2_1_2   ( clk , write2_29  , RELUout_F2_1_2  , Final_29_F2_1_2  );
OneRegister RAM_OUT_29_F2_2_1   ( clk , write2_29  , RELUout_F2_2_1  , Final_29_F2_2_1  );
OneRegister RAM_OUT_29_F2_2_2   ( clk , write2_29  , RELUout_F2_2_2  , Final_29_F2_2_2  );
OneRegister RAM_OUT_29_F3_1_1   ( clk , write2_29  , RELUout_F3_1_1  , Final_29_F3_1_1  );
OneRegister RAM_OUT_29_F3_1_2   ( clk , write2_29  , RELUout_F3_1_2  , Final_29_F3_1_2  );
OneRegister RAM_OUT_29_F3_2_1   ( clk , write2_29  , RELUout_F3_2_1  , Final_29_F3_2_1  );
OneRegister RAM_OUT_29_F3_2_2   ( clk , write2_29  , RELUout_F3_2_2  , Final_29_F3_2_2  );
OneRegister RAM_OUT_29_F4_1_1   ( clk , write2_29  , RELUout_F4_1_1  , Final_29_F4_1_1  );
OneRegister RAM_OUT_29_F4_1_2   ( clk , write2_29  , RELUout_F4_1_2  , Final_29_F4_1_2  );
OneRegister RAM_OUT_29_F4_2_1   ( clk , write2_29  , RELUout_F4_2_1  , Final_29_F4_2_1  );
OneRegister RAM_OUT_29_F4_2_2   ( clk , write2_29  , RELUout_F4_2_2  , Final_29_F4_2_2  );
OneRegister RAM_OUT_30_F1_1_1   ( clk , write2_30  , RELUout_F1_1_1  , Final_30_F1_1_1  );
OneRegister RAM_OUT_30_F1_1_2   ( clk , write2_30  , RELUout_F1_1_2  , Final_30_F1_1_2  );
OneRegister RAM_OUT_30_F1_2_1   ( clk , write2_30  , RELUout_F1_2_1  , Final_30_F1_2_1  );
OneRegister RAM_OUT_30_F1_2_2   ( clk , write2_30  , RELUout_F1_2_2  , Final_30_F1_2_2  );
OneRegister RAM_OUT_30_F2_1_1   ( clk , write2_30  , RELUout_F2_1_1  , Final_30_F2_1_1  );
OneRegister RAM_OUT_30_F2_1_2   ( clk , write2_30  , RELUout_F2_1_2  , Final_30_F2_1_2  );
OneRegister RAM_OUT_30_F2_2_1   ( clk , write2_30  , RELUout_F2_2_1  , Final_30_F2_2_1  );
OneRegister RAM_OUT_30_F2_2_2   ( clk , write2_30  , RELUout_F2_2_2  , Final_30_F2_2_2  );
OneRegister RAM_OUT_30_F3_1_1   ( clk , write2_30  , RELUout_F3_1_1  , Final_30_F3_1_1  );
OneRegister RAM_OUT_30_F3_1_2   ( clk , write2_30  , RELUout_F3_1_2  , Final_30_F3_1_2  );
OneRegister RAM_OUT_30_F3_2_1   ( clk , write2_30  , RELUout_F3_2_1  , Final_30_F3_2_1  );
OneRegister RAM_OUT_30_F3_2_2   ( clk , write2_30  , RELUout_F3_2_2  , Final_30_F3_2_2  );
OneRegister RAM_OUT_30_F4_1_1   ( clk , write2_30  , RELUout_F4_1_1  , Final_30_F4_1_1  );
OneRegister RAM_OUT_30_F4_1_2   ( clk , write2_30  , RELUout_F4_1_2  , Final_30_F4_1_2  );
OneRegister RAM_OUT_30_F4_2_1   ( clk , write2_30  , RELUout_F4_2_1  , Final_30_F4_2_1  );
OneRegister RAM_OUT_30_F4_2_2   ( clk , write2_30  , RELUout_F4_2_2  , Final_30_F4_2_2  );
OneRegister RAM_OUT_31_F1_1_1   ( clk , write2_31  , RELUout_F1_1_1  , Final_31_F1_1_1  );
OneRegister RAM_OUT_31_F1_1_2   ( clk , write2_31  , RELUout_F1_1_2  , Final_31_F1_1_2  );
OneRegister RAM_OUT_31_F1_2_1   ( clk , write2_31  , RELUout_F1_2_1  , Final_31_F1_2_1  );
OneRegister RAM_OUT_31_F1_2_2   ( clk , write2_31  , RELUout_F1_2_2  , Final_31_F1_2_2  );
OneRegister RAM_OUT_31_F2_1_1   ( clk , write2_31  , RELUout_F2_1_1  , Final_31_F2_1_1  );
OneRegister RAM_OUT_31_F2_1_2   ( clk , write2_31  , RELUout_F2_1_2  , Final_31_F2_1_2  );
OneRegister RAM_OUT_31_F2_2_1   ( clk , write2_31  , RELUout_F2_2_1  , Final_31_F2_2_1  );
OneRegister RAM_OUT_31_F2_2_2   ( clk , write2_31  , RELUout_F2_2_2  , Final_31_F2_2_2  );
OneRegister RAM_OUT_31_F3_1_1   ( clk , write2_31  , RELUout_F3_1_1  , Final_31_F3_1_1  );
OneRegister RAM_OUT_31_F3_1_2   ( clk , write2_31  , RELUout_F3_1_2  , Final_31_F3_1_2  );
OneRegister RAM_OUT_31_F3_2_1   ( clk , write2_31  , RELUout_F3_2_1  , Final_31_F3_2_1  );
OneRegister RAM_OUT_31_F3_2_2   ( clk , write2_31  , RELUout_F3_2_2  , Final_31_F3_2_2  );
OneRegister RAM_OUT_31_F4_1_1   ( clk , write2_31  , RELUout_F4_1_1  , Final_31_F4_1_1  );
OneRegister RAM_OUT_31_F4_1_2   ( clk , write2_31  , RELUout_F4_1_2  , Final_31_F4_1_2  );
OneRegister RAM_OUT_31_F4_2_1   ( clk , write2_31  , RELUout_F4_2_1  , Final_31_F4_2_1  );
OneRegister RAM_OUT_31_F4_2_2   ( clk , write2_31  , RELUout_F4_2_2  , Final_31_F4_2_2  );
OneRegister RAM_OUT_32_F1_1_1   ( clk , write2_32  , RELUout_F1_1_1  , Final_32_F1_1_1  );
OneRegister RAM_OUT_32_F1_1_2   ( clk , write2_32  , RELUout_F1_1_2  , Final_32_F1_1_2  );
OneRegister RAM_OUT_32_F1_2_1   ( clk , write2_32  , RELUout_F1_2_1  , Final_32_F1_2_1  );
OneRegister RAM_OUT_32_F1_2_2   ( clk , write2_32  , RELUout_F1_2_2  , Final_32_F1_2_2  );
OneRegister RAM_OUT_32_F2_1_1   ( clk , write2_32  , RELUout_F2_1_1  , Final_32_F2_1_1  );
OneRegister RAM_OUT_32_F2_1_2   ( clk , write2_32  , RELUout_F2_1_2  , Final_32_F2_1_2  );
OneRegister RAM_OUT_32_F2_2_1   ( clk , write2_32  , RELUout_F2_2_1  , Final_32_F2_2_1  );
OneRegister RAM_OUT_32_F2_2_2   ( clk , write2_32  , RELUout_F2_2_2  , Final_32_F2_2_2  );
OneRegister RAM_OUT_32_F3_1_1   ( clk , write2_32  , RELUout_F3_1_1  , Final_32_F3_1_1  );
OneRegister RAM_OUT_32_F3_1_2   ( clk , write2_32  , RELUout_F3_1_2  , Final_32_F3_1_2  );
OneRegister RAM_OUT_32_F3_2_1   ( clk , write2_32  , RELUout_F3_2_1  , Final_32_F3_2_1  );
OneRegister RAM_OUT_32_F3_2_2   ( clk , write2_32  , RELUout_F3_2_2  , Final_32_F3_2_2  );
OneRegister RAM_OUT_32_F4_1_1   ( clk , write2_32  , RELUout_F4_1_1  , Final_32_F4_1_1  );
OneRegister RAM_OUT_32_F4_1_2   ( clk , write2_32  , RELUout_F4_1_2  , Final_32_F4_1_2  );
OneRegister RAM_OUT_32_F4_2_1   ( clk , write2_32  , RELUout_F4_2_1  , Final_32_F4_2_1  );
OneRegister RAM_OUT_32_F4_2_2   ( clk , write2_32  , RELUout_F4_2_2  , Final_32_F4_2_2  );
OneRegister RAM_OUT_33_F1_1_1   ( clk , write2_33  , RELUout_F1_1_1  , Final_33_F1_1_1  );
OneRegister RAM_OUT_33_F1_1_2   ( clk , write2_33  , RELUout_F1_1_2  , Final_33_F1_1_2  );
OneRegister RAM_OUT_33_F1_2_1   ( clk , write2_33  , RELUout_F1_2_1  , Final_33_F1_2_1  );
OneRegister RAM_OUT_33_F1_2_2   ( clk , write2_33  , RELUout_F1_2_2  , Final_33_F1_2_2  );
OneRegister RAM_OUT_33_F2_1_1   ( clk , write2_33  , RELUout_F2_1_1  , Final_33_F2_1_1  );
OneRegister RAM_OUT_33_F2_1_2   ( clk , write2_33  , RELUout_F2_1_2  , Final_33_F2_1_2  );
OneRegister RAM_OUT_33_F2_2_1   ( clk , write2_33  , RELUout_F2_2_1  , Final_33_F2_2_1  );
OneRegister RAM_OUT_33_F2_2_2   ( clk , write2_33  , RELUout_F2_2_2  , Final_33_F2_2_2  );
OneRegister RAM_OUT_33_F3_1_1   ( clk , write2_33  , RELUout_F3_1_1  , Final_33_F3_1_1  );
OneRegister RAM_OUT_33_F3_1_2   ( clk , write2_33  , RELUout_F3_1_2  , Final_33_F3_1_2  );
OneRegister RAM_OUT_33_F3_2_1   ( clk , write2_33  , RELUout_F3_2_1  , Final_33_F3_2_1  );
OneRegister RAM_OUT_33_F3_2_2   ( clk , write2_33  , RELUout_F3_2_2  , Final_33_F3_2_2  );
OneRegister RAM_OUT_33_F4_1_1   ( clk , write2_33  , RELUout_F4_1_1  , Final_33_F4_1_1  );
OneRegister RAM_OUT_33_F4_1_2   ( clk , write2_33  , RELUout_F4_1_2  , Final_33_F4_1_2  );
OneRegister RAM_OUT_33_F4_2_1   ( clk , write2_33  , RELUout_F4_2_1  , Final_33_F4_2_1  );
OneRegister RAM_OUT_33_F4_2_2   ( clk , write2_33  , RELUout_F4_2_2  , Final_33_F4_2_2  );
OneRegister RAM_OUT_34_F1_1_1   ( clk , write2_34  , RELUout_F1_1_1  , Final_34_F1_1_1  );
OneRegister RAM_OUT_34_F1_1_2   ( clk , write2_34  , RELUout_F1_1_2  , Final_34_F1_1_2  );
OneRegister RAM_OUT_34_F1_2_1   ( clk , write2_34  , RELUout_F1_2_1  , Final_34_F1_2_1  );
OneRegister RAM_OUT_34_F1_2_2   ( clk , write2_34  , RELUout_F1_2_2  , Final_34_F1_2_2  );
OneRegister RAM_OUT_34_F2_1_1   ( clk , write2_34  , RELUout_F2_1_1  , Final_34_F2_1_1  );
OneRegister RAM_OUT_34_F2_1_2   ( clk , write2_34  , RELUout_F2_1_2  , Final_34_F2_1_2  );
OneRegister RAM_OUT_34_F2_2_1   ( clk , write2_34  , RELUout_F2_2_1  , Final_34_F2_2_1  );
OneRegister RAM_OUT_34_F2_2_2   ( clk , write2_34  , RELUout_F2_2_2  , Final_34_F2_2_2  );
OneRegister RAM_OUT_34_F3_1_1   ( clk , write2_34  , RELUout_F3_1_1  , Final_34_F3_1_1  );
OneRegister RAM_OUT_34_F3_1_2   ( clk , write2_34  , RELUout_F3_1_2  , Final_34_F3_1_2  );
OneRegister RAM_OUT_34_F3_2_1   ( clk , write2_34  , RELUout_F3_2_1  , Final_34_F3_2_1  );
OneRegister RAM_OUT_34_F3_2_2   ( clk , write2_34  , RELUout_F3_2_2  , Final_34_F3_2_2  );
OneRegister RAM_OUT_34_F4_1_1   ( clk , write2_34  , RELUout_F4_1_1  , Final_34_F4_1_1  );
OneRegister RAM_OUT_34_F4_1_2   ( clk , write2_34  , RELUout_F4_1_2  , Final_34_F4_1_2  );
OneRegister RAM_OUT_34_F4_2_1   ( clk , write2_34  , RELUout_F4_2_1  , Final_34_F4_2_1  );
OneRegister RAM_OUT_34_F4_2_2   ( clk , write2_34  , RELUout_F4_2_2  , Final_34_F4_2_2  );
OneRegister RAM_OUT_35_F1_1_1   ( clk , write2_35  , RELUout_F1_1_1  , Final_35_F1_1_1  );
OneRegister RAM_OUT_35_F1_1_2   ( clk , write2_35  , RELUout_F1_1_2  , Final_35_F1_1_2  );
OneRegister RAM_OUT_35_F1_2_1   ( clk , write2_35  , RELUout_F1_2_1  , Final_35_F1_2_1  );
OneRegister RAM_OUT_35_F1_2_2   ( clk , write2_35  , RELUout_F1_2_2  , Final_35_F1_2_2  );
OneRegister RAM_OUT_35_F2_1_1   ( clk , write2_35  , RELUout_F2_1_1  , Final_35_F2_1_1  );
OneRegister RAM_OUT_35_F2_1_2   ( clk , write2_35  , RELUout_F2_1_2  , Final_35_F2_1_2  );
OneRegister RAM_OUT_35_F2_2_1   ( clk , write2_35  , RELUout_F2_2_1  , Final_35_F2_2_1  );
OneRegister RAM_OUT_35_F2_2_2   ( clk , write2_35  , RELUout_F2_2_2  , Final_35_F2_2_2  );
OneRegister RAM_OUT_35_F3_1_1   ( clk , write2_35  , RELUout_F3_1_1  , Final_35_F3_1_1  );
OneRegister RAM_OUT_35_F3_1_2   ( clk , write2_35  , RELUout_F3_1_2  , Final_35_F3_1_2  );
OneRegister RAM_OUT_35_F3_2_1   ( clk , write2_35  , RELUout_F3_2_1  , Final_35_F3_2_1  );
OneRegister RAM_OUT_35_F3_2_2   ( clk , write2_35  , RELUout_F3_2_2  , Final_35_F3_2_2  );
OneRegister RAM_OUT_35_F4_1_1   ( clk , write2_35  , RELUout_F4_1_1  , Final_35_F4_1_1  );
OneRegister RAM_OUT_35_F4_1_2   ( clk , write2_35  , RELUout_F4_1_2  , Final_35_F4_1_2  );
OneRegister RAM_OUT_35_F4_2_1   ( clk , write2_35  , RELUout_F4_2_1  , Final_35_F4_2_1  );
OneRegister RAM_OUT_35_F4_2_2   ( clk , write2_35  , RELUout_F4_2_2  , Final_35_F4_2_2  );
OneRegister RAM_OUT_36_F1_1_1   ( clk , write2_36  , RELUout_F1_1_1  , Final_36_F1_1_1  );
OneRegister RAM_OUT_36_F1_1_2   ( clk , write2_36  , RELUout_F1_1_2  , Final_36_F1_1_2  );
OneRegister RAM_OUT_36_F1_2_1   ( clk , write2_36  , RELUout_F1_2_1  , Final_36_F1_2_1  );
OneRegister RAM_OUT_36_F1_2_2   ( clk , write2_36  , RELUout_F1_2_2  , Final_36_F1_2_2  );
OneRegister RAM_OUT_36_F2_1_1   ( clk , write2_36  , RELUout_F2_1_1  , Final_36_F2_1_1  );
OneRegister RAM_OUT_36_F2_1_2   ( clk , write2_36  , RELUout_F2_1_2  , Final_36_F2_1_2  );
OneRegister RAM_OUT_36_F2_2_1   ( clk , write2_36  , RELUout_F2_2_1  , Final_36_F2_2_1  );
OneRegister RAM_OUT_36_F2_2_2   ( clk , write2_36  , RELUout_F2_2_2  , Final_36_F2_2_2  );
OneRegister RAM_OUT_36_F3_1_1   ( clk , write2_36  , RELUout_F3_1_1  , Final_36_F3_1_1  );
OneRegister RAM_OUT_36_F3_1_2   ( clk , write2_36  , RELUout_F3_1_2  , Final_36_F3_1_2  );
OneRegister RAM_OUT_36_F3_2_1   ( clk , write2_36  , RELUout_F3_2_1  , Final_36_F3_2_1  );
OneRegister RAM_OUT_36_F3_2_2   ( clk , write2_36  , RELUout_F3_2_2  , Final_36_F3_2_2  );
OneRegister RAM_OUT_36_F4_1_1   ( clk , write2_36  , RELUout_F4_1_1  , Final_36_F4_1_1  );
OneRegister RAM_OUT_36_F4_1_2   ( clk , write2_36  , RELUout_F4_1_2  , Final_36_F4_1_2  );
OneRegister RAM_OUT_36_F4_2_1   ( clk , write2_36  , RELUout_F4_2_1  , Final_36_F4_2_1  );
OneRegister RAM_OUT_36_F4_2_2   ( clk , write2_36  , RELUout_F4_2_2  , Final_36_F4_2_2  );
OneRegister RAM_OUT_37_F1_1_1   ( clk , write2_37  , RELUout_F1_1_1  , Final_37_F1_1_1  );
OneRegister RAM_OUT_37_F1_1_2   ( clk , write2_37  , RELUout_F1_1_2  , Final_37_F1_1_2  );
OneRegister RAM_OUT_37_F1_2_1   ( clk , write2_37  , RELUout_F1_2_1  , Final_37_F1_2_1  );
OneRegister RAM_OUT_37_F1_2_2   ( clk , write2_37  , RELUout_F1_2_2  , Final_37_F1_2_2  );
OneRegister RAM_OUT_37_F2_1_1   ( clk , write2_37  , RELUout_F2_1_1  , Final_37_F2_1_1  );
OneRegister RAM_OUT_37_F2_1_2   ( clk , write2_37  , RELUout_F2_1_2  , Final_37_F2_1_2  );
OneRegister RAM_OUT_37_F2_2_1   ( clk , write2_37  , RELUout_F2_2_1  , Final_37_F2_2_1  );
OneRegister RAM_OUT_37_F2_2_2   ( clk , write2_37  , RELUout_F2_2_2  , Final_37_F2_2_2  );
OneRegister RAM_OUT_37_F3_1_1   ( clk , write2_37  , RELUout_F3_1_1  , Final_37_F3_1_1  );
OneRegister RAM_OUT_37_F3_1_2   ( clk , write2_37  , RELUout_F3_1_2  , Final_37_F3_1_2  );
OneRegister RAM_OUT_37_F3_2_1   ( clk , write2_37  , RELUout_F3_2_1  , Final_37_F3_2_1  );
OneRegister RAM_OUT_37_F3_2_2   ( clk , write2_37  , RELUout_F3_2_2  , Final_37_F3_2_2  );
OneRegister RAM_OUT_37_F4_1_1   ( clk , write2_37  , RELUout_F4_1_1  , Final_37_F4_1_1  );
OneRegister RAM_OUT_37_F4_1_2   ( clk , write2_37  , RELUout_F4_1_2  , Final_37_F4_1_2  );
OneRegister RAM_OUT_37_F4_2_1   ( clk , write2_37  , RELUout_F4_2_1  , Final_37_F4_2_1  );
OneRegister RAM_OUT_37_F4_2_2   ( clk , write2_37  , RELUout_F4_2_2  , Final_37_F4_2_2  );
OneRegister RAM_OUT_38_F1_1_1   ( clk , write2_38  , RELUout_F1_1_1  , Final_38_F1_1_1  );
OneRegister RAM_OUT_38_F1_1_2   ( clk , write2_38  , RELUout_F1_1_2  , Final_38_F1_1_2  );
OneRegister RAM_OUT_38_F1_2_1   ( clk , write2_38  , RELUout_F1_2_1  , Final_38_F1_2_1  );
OneRegister RAM_OUT_38_F1_2_2   ( clk , write2_38  , RELUout_F1_2_2  , Final_38_F1_2_2  );
OneRegister RAM_OUT_38_F2_1_1   ( clk , write2_38  , RELUout_F2_1_1  , Final_38_F2_1_1  );
OneRegister RAM_OUT_38_F2_1_2   ( clk , write2_38  , RELUout_F2_1_2  , Final_38_F2_1_2  );
OneRegister RAM_OUT_38_F2_2_1   ( clk , write2_38  , RELUout_F2_2_1  , Final_38_F2_2_1  );
OneRegister RAM_OUT_38_F2_2_2   ( clk , write2_38  , RELUout_F2_2_2  , Final_38_F2_2_2  );
OneRegister RAM_OUT_38_F3_1_1   ( clk , write2_38  , RELUout_F3_1_1  , Final_38_F3_1_1  );
OneRegister RAM_OUT_38_F3_1_2   ( clk , write2_38  , RELUout_F3_1_2  , Final_38_F3_1_2  );
OneRegister RAM_OUT_38_F3_2_1   ( clk , write2_38  , RELUout_F3_2_1  , Final_38_F3_2_1  );
OneRegister RAM_OUT_38_F3_2_2   ( clk , write2_38  , RELUout_F3_2_2  , Final_38_F3_2_2  );
OneRegister RAM_OUT_38_F4_1_1   ( clk , write2_38  , RELUout_F4_1_1  , Final_38_F4_1_1  );
OneRegister RAM_OUT_38_F4_1_2   ( clk , write2_38  , RELUout_F4_1_2  , Final_38_F4_1_2  );
OneRegister RAM_OUT_38_F4_2_1   ( clk , write2_38  , RELUout_F4_2_1  , Final_38_F4_2_1  );
OneRegister RAM_OUT_38_F4_2_2   ( clk , write2_38  , RELUout_F4_2_2  , Final_38_F4_2_2  );
OneRegister RAM_OUT_39_F1_1_1   ( clk , write2_39  , RELUout_F1_1_1  , Final_39_F1_1_1  );
OneRegister RAM_OUT_39_F1_1_2   ( clk , write2_39  , RELUout_F1_1_2  , Final_39_F1_1_2  );
OneRegister RAM_OUT_39_F1_2_1   ( clk , write2_39  , RELUout_F1_2_1  , Final_39_F1_2_1  );
OneRegister RAM_OUT_39_F1_2_2   ( clk , write2_39  , RELUout_F1_2_2  , Final_39_F1_2_2  );
OneRegister RAM_OUT_39_F2_1_1   ( clk , write2_39  , RELUout_F2_1_1  , Final_39_F2_1_1  );
OneRegister RAM_OUT_39_F2_1_2   ( clk , write2_39  , RELUout_F2_1_2  , Final_39_F2_1_2  );
OneRegister RAM_OUT_39_F2_2_1   ( clk , write2_39  , RELUout_F2_2_1  , Final_39_F2_2_1  );
OneRegister RAM_OUT_39_F2_2_2   ( clk , write2_39  , RELUout_F2_2_2  , Final_39_F2_2_2  );
OneRegister RAM_OUT_39_F3_1_1   ( clk , write2_39  , RELUout_F3_1_1  , Final_39_F3_1_1  );
OneRegister RAM_OUT_39_F3_1_2   ( clk , write2_39  , RELUout_F3_1_2  , Final_39_F3_1_2  );
OneRegister RAM_OUT_39_F3_2_1   ( clk , write2_39  , RELUout_F3_2_1  , Final_39_F3_2_1  );
OneRegister RAM_OUT_39_F3_2_2   ( clk , write2_39  , RELUout_F3_2_2  , Final_39_F3_2_2  );
OneRegister RAM_OUT_39_F4_1_1   ( clk , write2_39  , RELUout_F4_1_1  , Final_39_F4_1_1  );
OneRegister RAM_OUT_39_F4_1_2   ( clk , write2_39  , RELUout_F4_1_2  , Final_39_F4_1_2  );
OneRegister RAM_OUT_39_F4_2_1   ( clk , write2_39  , RELUout_F4_2_1  , Final_39_F4_2_1  );
OneRegister RAM_OUT_39_F4_2_2   ( clk , write2_39  , RELUout_F4_2_2  , Final_39_F4_2_2  );
OneRegister RAM_OUT_40_F1_1_1   ( clk , write2_40  , RELUout_F1_1_1  , Final_40_F1_1_1  );
OneRegister RAM_OUT_40_F1_1_2   ( clk , write2_40  , RELUout_F1_1_2  , Final_40_F1_1_2  );
OneRegister RAM_OUT_40_F1_2_1   ( clk , write2_40  , RELUout_F1_2_1  , Final_40_F1_2_1  );
OneRegister RAM_OUT_40_F1_2_2   ( clk , write2_40  , RELUout_F1_2_2  , Final_40_F1_2_2  );
OneRegister RAM_OUT_40_F2_1_1   ( clk , write2_40  , RELUout_F2_1_1  , Final_40_F2_1_1  );
OneRegister RAM_OUT_40_F2_1_2   ( clk , write2_40  , RELUout_F2_1_2  , Final_40_F2_1_2  );
OneRegister RAM_OUT_40_F2_2_1   ( clk , write2_40  , RELUout_F2_2_1  , Final_40_F2_2_1  );
OneRegister RAM_OUT_40_F2_2_2   ( clk , write2_40  , RELUout_F2_2_2  , Final_40_F2_2_2  );
OneRegister RAM_OUT_40_F3_1_1   ( clk , write2_40  , RELUout_F3_1_1  , Final_40_F3_1_1  );
OneRegister RAM_OUT_40_F3_1_2   ( clk , write2_40  , RELUout_F3_1_2  , Final_40_F3_1_2  );
OneRegister RAM_OUT_40_F3_2_1   ( clk , write2_40  , RELUout_F3_2_1  , Final_40_F3_2_1  );
OneRegister RAM_OUT_40_F3_2_2   ( clk , write2_40  , RELUout_F3_2_2  , Final_40_F3_2_2  );
OneRegister RAM_OUT_40_F4_1_1   ( clk , write2_40  , RELUout_F4_1_1  , Final_40_F4_1_1  );
OneRegister RAM_OUT_40_F4_1_2   ( clk , write2_40  , RELUout_F4_1_2  , Final_40_F4_1_2  );
OneRegister RAM_OUT_40_F4_2_1   ( clk , write2_40  , RELUout_F4_2_1  , Final_40_F4_2_1  );
OneRegister RAM_OUT_40_F4_2_2   ( clk , write2_40  , RELUout_F4_2_2  , Final_40_F4_2_2  );
OneRegister RAM_OUT_41_F1_1_1   ( clk , write2_41  , RELUout_F1_1_1  , Final_41_F1_1_1  );
OneRegister RAM_OUT_41_F1_1_2   ( clk , write2_41  , RELUout_F1_1_2  , Final_41_F1_1_2  );
OneRegister RAM_OUT_41_F1_2_1   ( clk , write2_41  , RELUout_F1_2_1  , Final_41_F1_2_1  );
OneRegister RAM_OUT_41_F1_2_2   ( clk , write2_41  , RELUout_F1_2_2  , Final_41_F1_2_2  );
OneRegister RAM_OUT_41_F2_1_1   ( clk , write2_41  , RELUout_F2_1_1  , Final_41_F2_1_1  );
OneRegister RAM_OUT_41_F2_1_2   ( clk , write2_41  , RELUout_F2_1_2  , Final_41_F2_1_2  );
OneRegister RAM_OUT_41_F2_2_1   ( clk , write2_41  , RELUout_F2_2_1  , Final_41_F2_2_1  );
OneRegister RAM_OUT_41_F2_2_2   ( clk , write2_41  , RELUout_F2_2_2  , Final_41_F2_2_2  );
OneRegister RAM_OUT_41_F3_1_1   ( clk , write2_41  , RELUout_F3_1_1  , Final_41_F3_1_1  );
OneRegister RAM_OUT_41_F3_1_2   ( clk , write2_41  , RELUout_F3_1_2  , Final_41_F3_1_2  );
OneRegister RAM_OUT_41_F3_2_1   ( clk , write2_41  , RELUout_F3_2_1  , Final_41_F3_2_1  );
OneRegister RAM_OUT_41_F3_2_2   ( clk , write2_41  , RELUout_F3_2_2  , Final_41_F3_2_2  );
OneRegister RAM_OUT_41_F4_1_1   ( clk , write2_41  , RELUout_F4_1_1  , Final_41_F4_1_1  );
OneRegister RAM_OUT_41_F4_1_2   ( clk , write2_41  , RELUout_F4_1_2  , Final_41_F4_1_2  );
OneRegister RAM_OUT_41_F4_2_1   ( clk , write2_41  , RELUout_F4_2_1  , Final_41_F4_2_1  );
OneRegister RAM_OUT_41_F4_2_2   ( clk , write2_41  , RELUout_F4_2_2  , Final_41_F4_2_2  );
OneRegister RAM_OUT_42_F1_1_1   ( clk , write2_42  , RELUout_F1_1_1  , Final_42_F1_1_1  );
OneRegister RAM_OUT_42_F1_1_2   ( clk , write2_42  , RELUout_F1_1_2  , Final_42_F1_1_2  );
OneRegister RAM_OUT_42_F1_2_1   ( clk , write2_42  , RELUout_F1_2_1  , Final_42_F1_2_1  );
OneRegister RAM_OUT_42_F1_2_2   ( clk , write2_42  , RELUout_F1_2_2  , Final_42_F1_2_2  );
OneRegister RAM_OUT_42_F2_1_1   ( clk , write2_42  , RELUout_F2_1_1  , Final_42_F2_1_1  );
OneRegister RAM_OUT_42_F2_1_2   ( clk , write2_42  , RELUout_F2_1_2  , Final_42_F2_1_2  );
OneRegister RAM_OUT_42_F2_2_1   ( clk , write2_42  , RELUout_F2_2_1  , Final_42_F2_2_1  );
OneRegister RAM_OUT_42_F2_2_2   ( clk , write2_42  , RELUout_F2_2_2  , Final_42_F2_2_2  );
OneRegister RAM_OUT_42_F3_1_1   ( clk , write2_42  , RELUout_F3_1_1  , Final_42_F3_1_1  );
OneRegister RAM_OUT_42_F3_1_2   ( clk , write2_42  , RELUout_F3_1_2  , Final_42_F3_1_2  );
OneRegister RAM_OUT_42_F3_2_1   ( clk , write2_42  , RELUout_F3_2_1  , Final_42_F3_2_1  );
OneRegister RAM_OUT_42_F3_2_2   ( clk , write2_42  , RELUout_F3_2_2  , Final_42_F3_2_2  );
OneRegister RAM_OUT_42_F4_1_1   ( clk , write2_42  , RELUout_F4_1_1  , Final_42_F4_1_1  );
OneRegister RAM_OUT_42_F4_1_2   ( clk , write2_42  , RELUout_F4_1_2  , Final_42_F4_1_2  );
OneRegister RAM_OUT_42_F4_2_1   ( clk , write2_42  , RELUout_F4_2_1  , Final_42_F4_2_1  );
OneRegister RAM_OUT_42_F4_2_2   ( clk , write2_42  , RELUout_F4_2_2  , Final_42_F4_2_2  );
OneRegister RAM_OUT_43_F1_1_1   ( clk , write2_43  , RELUout_F1_1_1  , Final_43_F1_1_1  );
OneRegister RAM_OUT_43_F1_1_2   ( clk , write2_43  , RELUout_F1_1_2  , Final_43_F1_1_2  );
OneRegister RAM_OUT_43_F1_2_1   ( clk , write2_43  , RELUout_F1_2_1  , Final_43_F1_2_1  );
OneRegister RAM_OUT_43_F1_2_2   ( clk , write2_43  , RELUout_F1_2_2  , Final_43_F1_2_2  );
OneRegister RAM_OUT_43_F2_1_1   ( clk , write2_43  , RELUout_F2_1_1  , Final_43_F2_1_1  );
OneRegister RAM_OUT_43_F2_1_2   ( clk , write2_43  , RELUout_F2_1_2  , Final_43_F2_1_2  );
OneRegister RAM_OUT_43_F2_2_1   ( clk , write2_43  , RELUout_F2_2_1  , Final_43_F2_2_1  );
OneRegister RAM_OUT_43_F2_2_2   ( clk , write2_43  , RELUout_F2_2_2  , Final_43_F2_2_2  );
OneRegister RAM_OUT_43_F3_1_1   ( clk , write2_43  , RELUout_F3_1_1  , Final_43_F3_1_1  );
OneRegister RAM_OUT_43_F3_1_2   ( clk , write2_43  , RELUout_F3_1_2  , Final_43_F3_1_2  );
OneRegister RAM_OUT_43_F3_2_1   ( clk , write2_43  , RELUout_F3_2_1  , Final_43_F3_2_1  );
OneRegister RAM_OUT_43_F3_2_2   ( clk , write2_43  , RELUout_F3_2_2  , Final_43_F3_2_2  );
OneRegister RAM_OUT_43_F4_1_1   ( clk , write2_43  , RELUout_F4_1_1  , Final_43_F4_1_1  );
OneRegister RAM_OUT_43_F4_1_2   ( clk , write2_43  , RELUout_F4_1_2  , Final_43_F4_1_2  );
OneRegister RAM_OUT_43_F4_2_1   ( clk , write2_43  , RELUout_F4_2_1  , Final_43_F4_2_1  );
OneRegister RAM_OUT_43_F4_2_2   ( clk , write2_43  , RELUout_F4_2_2  , Final_43_F4_2_2  );
OneRegister RAM_OUT_44_F1_1_1   ( clk , write2_44  , RELUout_F1_1_1  , Final_44_F1_1_1  );
OneRegister RAM_OUT_44_F1_1_2   ( clk , write2_44  , RELUout_F1_1_2  , Final_44_F1_1_2  );
OneRegister RAM_OUT_44_F1_2_1   ( clk , write2_44  , RELUout_F1_2_1  , Final_44_F1_2_1  );
OneRegister RAM_OUT_44_F1_2_2   ( clk , write2_44  , RELUout_F1_2_2  , Final_44_F1_2_2  );
OneRegister RAM_OUT_44_F2_1_1   ( clk , write2_44  , RELUout_F2_1_1  , Final_44_F2_1_1  );
OneRegister RAM_OUT_44_F2_1_2   ( clk , write2_44  , RELUout_F2_1_2  , Final_44_F2_1_2  );
OneRegister RAM_OUT_44_F2_2_1   ( clk , write2_44  , RELUout_F2_2_1  , Final_44_F2_2_1  );
OneRegister RAM_OUT_44_F2_2_2   ( clk , write2_44  , RELUout_F2_2_2  , Final_44_F2_2_2  );
OneRegister RAM_OUT_44_F3_1_1   ( clk , write2_44  , RELUout_F3_1_1  , Final_44_F3_1_1  );
OneRegister RAM_OUT_44_F3_1_2   ( clk , write2_44  , RELUout_F3_1_2  , Final_44_F3_1_2  );
OneRegister RAM_OUT_44_F3_2_1   ( clk , write2_44  , RELUout_F3_2_1  , Final_44_F3_2_1  );
OneRegister RAM_OUT_44_F3_2_2   ( clk , write2_44  , RELUout_F3_2_2  , Final_44_F3_2_2  );
OneRegister RAM_OUT_44_F4_1_1   ( clk , write2_44  , RELUout_F4_1_1  , Final_44_F4_1_1  );
OneRegister RAM_OUT_44_F4_1_2   ( clk , write2_44  , RELUout_F4_1_2  , Final_44_F4_1_2  );
OneRegister RAM_OUT_44_F4_2_1   ( clk , write2_44  , RELUout_F4_2_1  , Final_44_F4_2_1  );
OneRegister RAM_OUT_44_F4_2_2   ( clk , write2_44  , RELUout_F4_2_2  , Final_44_F4_2_2  );
OneRegister RAM_OUT_45_F1_1_1   ( clk , write2_45  , RELUout_F1_1_1  , Final_45_F1_1_1  );
OneRegister RAM_OUT_45_F1_1_2   ( clk , write2_45  , RELUout_F1_1_2  , Final_45_F1_1_2  );
OneRegister RAM_OUT_45_F1_2_1   ( clk , write2_45  , RELUout_F1_2_1  , Final_45_F1_2_1  );
OneRegister RAM_OUT_45_F1_2_2   ( clk , write2_45  , RELUout_F1_2_2  , Final_45_F1_2_2  );
OneRegister RAM_OUT_45_F2_1_1   ( clk , write2_45  , RELUout_F2_1_1  , Final_45_F2_1_1  );
OneRegister RAM_OUT_45_F2_1_2   ( clk , write2_45  , RELUout_F2_1_2  , Final_45_F2_1_2  );
OneRegister RAM_OUT_45_F2_2_1   ( clk , write2_45  , RELUout_F2_2_1  , Final_45_F2_2_1  );
OneRegister RAM_OUT_45_F2_2_2   ( clk , write2_45  , RELUout_F2_2_2  , Final_45_F2_2_2  );
OneRegister RAM_OUT_45_F3_1_1   ( clk , write2_45  , RELUout_F3_1_1  , Final_45_F3_1_1  );
OneRegister RAM_OUT_45_F3_1_2   ( clk , write2_45  , RELUout_F3_1_2  , Final_45_F3_1_2  );
OneRegister RAM_OUT_45_F3_2_1   ( clk , write2_45  , RELUout_F3_2_1  , Final_45_F3_2_1  );
OneRegister RAM_OUT_45_F3_2_2   ( clk , write2_45  , RELUout_F3_2_2  , Final_45_F3_2_2  );
OneRegister RAM_OUT_45_F4_1_1   ( clk , write2_45  , RELUout_F4_1_1  , Final_45_F4_1_1  );
OneRegister RAM_OUT_45_F4_1_2   ( clk , write2_45  , RELUout_F4_1_2  , Final_45_F4_1_2  );
OneRegister RAM_OUT_45_F4_2_1   ( clk , write2_45  , RELUout_F4_2_1  , Final_45_F4_2_1  );
OneRegister RAM_OUT_45_F4_2_2   ( clk , write2_45  , RELUout_F4_2_2  , Final_45_F4_2_2  );
OneRegister RAM_OUT_46_F1_1_1   ( clk , write2_46  , RELUout_F1_1_1  , Final_46_F1_1_1  );
OneRegister RAM_OUT_46_F1_1_2   ( clk , write2_46  , RELUout_F1_1_2  , Final_46_F1_1_2  );
OneRegister RAM_OUT_46_F1_2_1   ( clk , write2_46  , RELUout_F1_2_1  , Final_46_F1_2_1  );
OneRegister RAM_OUT_46_F1_2_2   ( clk , write2_46  , RELUout_F1_2_2  , Final_46_F1_2_2  );
OneRegister RAM_OUT_46_F2_1_1   ( clk , write2_46  , RELUout_F2_1_1  , Final_46_F2_1_1  );
OneRegister RAM_OUT_46_F2_1_2   ( clk , write2_46  , RELUout_F2_1_2  , Final_46_F2_1_2  );
OneRegister RAM_OUT_46_F2_2_1   ( clk , write2_46  , RELUout_F2_2_1  , Final_46_F2_2_1  );
OneRegister RAM_OUT_46_F2_2_2   ( clk , write2_46  , RELUout_F2_2_2  , Final_46_F2_2_2  );
OneRegister RAM_OUT_46_F3_1_1   ( clk , write2_46  , RELUout_F3_1_1  , Final_46_F3_1_1  );
OneRegister RAM_OUT_46_F3_1_2   ( clk , write2_46  , RELUout_F3_1_2  , Final_46_F3_1_2  );
OneRegister RAM_OUT_46_F3_2_1   ( clk , write2_46  , RELUout_F3_2_1  , Final_46_F3_2_1  );
OneRegister RAM_OUT_46_F3_2_2   ( clk , write2_46  , RELUout_F3_2_2  , Final_46_F3_2_2  );
OneRegister RAM_OUT_46_F4_1_1   ( clk , write2_46  , RELUout_F4_1_1  , Final_46_F4_1_1  );
OneRegister RAM_OUT_46_F4_1_2   ( clk , write2_46  , RELUout_F4_1_2  , Final_46_F4_1_2  );
OneRegister RAM_OUT_46_F4_2_1   ( clk , write2_46  , RELUout_F4_2_1  , Final_46_F4_2_1  );
OneRegister RAM_OUT_46_F4_2_2   ( clk , write2_46  , RELUout_F4_2_2  , Final_46_F4_2_2  );
OneRegister RAM_OUT_47_F1_1_1   ( clk , write2_47  , RELUout_F1_1_1  , Final_47_F1_1_1  );
OneRegister RAM_OUT_47_F1_1_2   ( clk , write2_47  , RELUout_F1_1_2  , Final_47_F1_1_2  );
OneRegister RAM_OUT_47_F1_2_1   ( clk , write2_47  , RELUout_F1_2_1  , Final_47_F1_2_1  );
OneRegister RAM_OUT_47_F1_2_2   ( clk , write2_47  , RELUout_F1_2_2  , Final_47_F1_2_2  );
OneRegister RAM_OUT_47_F2_1_1   ( clk , write2_47  , RELUout_F2_1_1  , Final_47_F2_1_1  );
OneRegister RAM_OUT_47_F2_1_2   ( clk , write2_47  , RELUout_F2_1_2  , Final_47_F2_1_2  );
OneRegister RAM_OUT_47_F2_2_1   ( clk , write2_47  , RELUout_F2_2_1  , Final_47_F2_2_1  );
OneRegister RAM_OUT_47_F2_2_2   ( clk , write2_47  , RELUout_F2_2_2  , Final_47_F2_2_2  );
OneRegister RAM_OUT_47_F3_1_1   ( clk , write2_47  , RELUout_F3_1_1  , Final_47_F3_1_1  );
OneRegister RAM_OUT_47_F3_1_2   ( clk , write2_47  , RELUout_F3_1_2  , Final_47_F3_1_2  );
OneRegister RAM_OUT_47_F3_2_1   ( clk , write2_47  , RELUout_F3_2_1  , Final_47_F3_2_1  );
OneRegister RAM_OUT_47_F3_2_2   ( clk , write2_47  , RELUout_F3_2_2  , Final_47_F3_2_2  );
OneRegister RAM_OUT_47_F4_1_1   ( clk , write2_47  , RELUout_F4_1_1  , Final_47_F4_1_1  );
OneRegister RAM_OUT_47_F4_1_2   ( clk , write2_47  , RELUout_F4_1_2  , Final_47_F4_1_2  );
OneRegister RAM_OUT_47_F4_2_1   ( clk , write2_47  , RELUout_F4_2_1  , Final_47_F4_2_1  );
OneRegister RAM_OUT_47_F4_2_2   ( clk , write2_47  , RELUout_F4_2_2  , Final_47_F4_2_2  );
OneRegister RAM_OUT_48_F1_1_1   ( clk , write2_48  , RELUout_F1_1_1  , Final_48_F1_1_1  );
OneRegister RAM_OUT_48_F1_1_2   ( clk , write2_48  , RELUout_F1_1_2  , Final_48_F1_1_2  );
OneRegister RAM_OUT_48_F1_2_1   ( clk , write2_48  , RELUout_F1_2_1  , Final_48_F1_2_1  );
OneRegister RAM_OUT_48_F1_2_2   ( clk , write2_48  , RELUout_F1_2_2  , Final_48_F1_2_2  );
OneRegister RAM_OUT_48_F2_1_1   ( clk , write2_48  , RELUout_F2_1_1  , Final_48_F2_1_1  );
OneRegister RAM_OUT_48_F2_1_2   ( clk , write2_48  , RELUout_F2_1_2  , Final_48_F2_1_2  );
OneRegister RAM_OUT_48_F2_2_1   ( clk , write2_48  , RELUout_F2_2_1  , Final_48_F2_2_1  );
OneRegister RAM_OUT_48_F2_2_2   ( clk , write2_48  , RELUout_F2_2_2  , Final_48_F2_2_2  );
OneRegister RAM_OUT_48_F3_1_1   ( clk , write2_48  , RELUout_F3_1_1  , Final_48_F3_1_1  );
OneRegister RAM_OUT_48_F3_1_2   ( clk , write2_48  , RELUout_F3_1_2  , Final_48_F3_1_2  );
OneRegister RAM_OUT_48_F3_2_1   ( clk , write2_48  , RELUout_F3_2_1  , Final_48_F3_2_1  );
OneRegister RAM_OUT_48_F3_2_2   ( clk , write2_48  , RELUout_F3_2_2  , Final_48_F3_2_2  );
OneRegister RAM_OUT_48_F4_1_1   ( clk , write2_48  , RELUout_F4_1_1  , Final_48_F4_1_1  );
OneRegister RAM_OUT_48_F4_1_2   ( clk , write2_48  , RELUout_F4_1_2  , Final_48_F4_1_2  );
OneRegister RAM_OUT_48_F4_2_1   ( clk , write2_48  , RELUout_F4_2_1  , Final_48_F4_2_1  );
OneRegister RAM_OUT_48_F4_2_2   ( clk , write2_48  , RELUout_F4_2_2  , Final_48_F4_2_2  );
OneRegister RAM_OUT_49_F1_1_1   ( clk , write2_49  , RELUout_F1_1_1  , Final_49_F1_1_1  );
OneRegister RAM_OUT_49_F1_1_2   ( clk , write2_49  , RELUout_F1_1_2  , Final_49_F1_1_2  );
OneRegister RAM_OUT_49_F1_2_1   ( clk , write2_49  , RELUout_F1_2_1  , Final_49_F1_2_1  );
OneRegister RAM_OUT_49_F1_2_2   ( clk , write2_49  , RELUout_F1_2_2  , Final_49_F1_2_2  );
OneRegister RAM_OUT_49_F2_1_1   ( clk , write2_49  , RELUout_F2_1_1  , Final_49_F2_1_1  );
OneRegister RAM_OUT_49_F2_1_2   ( clk , write2_49  , RELUout_F2_1_2  , Final_49_F2_1_2  );
OneRegister RAM_OUT_49_F2_2_1   ( clk , write2_49  , RELUout_F2_2_1  , Final_49_F2_2_1  );
OneRegister RAM_OUT_49_F2_2_2   ( clk , write2_49  , RELUout_F2_2_2  , Final_49_F2_2_2  );
OneRegister RAM_OUT_49_F3_1_1   ( clk , write2_49  , RELUout_F3_1_1  , Final_49_F3_1_1  );
OneRegister RAM_OUT_49_F3_1_2   ( clk , write2_49  , RELUout_F3_1_2  , Final_49_F3_1_2  );
OneRegister RAM_OUT_49_F3_2_1   ( clk , write2_49  , RELUout_F3_2_1  , Final_49_F3_2_1  );
OneRegister RAM_OUT_49_F3_2_2   ( clk , write2_49  , RELUout_F3_2_2  , Final_49_F3_2_2  );
OneRegister RAM_OUT_49_F4_1_1   ( clk , write2_49  , RELUout_F4_1_1  , Final_49_F4_1_1  );
OneRegister RAM_OUT_49_F4_1_2   ( clk , write2_49  , RELUout_F4_1_2  , Final_49_F4_1_2  );
OneRegister RAM_OUT_49_F4_2_1   ( clk , write2_49  , RELUout_F4_2_1  , Final_49_F4_2_1  );
OneRegister RAM_OUT_49_F4_2_2   ( clk , write2_49  , RELUout_F4_2_2  , Final_49_F4_2_2  );
OneRegister RAM_OUT_50_F1_1_1   ( clk , write2_50  , RELUout_F1_1_1  , Final_50_F1_1_1  );
OneRegister RAM_OUT_50_F1_1_2   ( clk , write2_50  , RELUout_F1_1_2  , Final_50_F1_1_2  );
OneRegister RAM_OUT_50_F1_2_1   ( clk , write2_50  , RELUout_F1_2_1  , Final_50_F1_2_1  );
OneRegister RAM_OUT_50_F1_2_2   ( clk , write2_50  , RELUout_F1_2_2  , Final_50_F1_2_2  );
OneRegister RAM_OUT_50_F2_1_1   ( clk , write2_50  , RELUout_F2_1_1  , Final_50_F2_1_1  );
OneRegister RAM_OUT_50_F2_1_2   ( clk , write2_50  , RELUout_F2_1_2  , Final_50_F2_1_2  );
OneRegister RAM_OUT_50_F2_2_1   ( clk , write2_50  , RELUout_F2_2_1  , Final_50_F2_2_1  );
OneRegister RAM_OUT_50_F2_2_2   ( clk , write2_50  , RELUout_F2_2_2  , Final_50_F2_2_2  );
OneRegister RAM_OUT_50_F3_1_1   ( clk , write2_50  , RELUout_F3_1_1  , Final_50_F3_1_1  );
OneRegister RAM_OUT_50_F3_1_2   ( clk , write2_50  , RELUout_F3_1_2  , Final_50_F3_1_2  );
OneRegister RAM_OUT_50_F3_2_1   ( clk , write2_50  , RELUout_F3_2_1  , Final_50_F3_2_1  );
OneRegister RAM_OUT_50_F3_2_2   ( clk , write2_50  , RELUout_F3_2_2  , Final_50_F3_2_2  );
OneRegister RAM_OUT_50_F4_1_1   ( clk , write2_50  , RELUout_F4_1_1  , Final_50_F4_1_1  );
OneRegister RAM_OUT_50_F4_1_2   ( clk , write2_50  , RELUout_F4_1_2  , Final_50_F4_1_2  );
OneRegister RAM_OUT_50_F4_2_1   ( clk , write2_50  , RELUout_F4_2_1  , Final_50_F4_2_1  );
OneRegister RAM_OUT_50_F4_2_2   ( clk , write2_50  , RELUout_F4_2_2  , Final_50_F4_2_2  );
OneRegister RAM_OUT_51_F1_1_1   ( clk , write2_51  , RELUout_F1_1_1  , Final_51_F1_1_1  );
OneRegister RAM_OUT_51_F1_1_2   ( clk , write2_51  , RELUout_F1_1_2  , Final_51_F1_1_2  );
OneRegister RAM_OUT_51_F1_2_1   ( clk , write2_51  , RELUout_F1_2_1  , Final_51_F1_2_1  );
OneRegister RAM_OUT_51_F1_2_2   ( clk , write2_51  , RELUout_F1_2_2  , Final_51_F1_2_2  );
OneRegister RAM_OUT_51_F2_1_1   ( clk , write2_51  , RELUout_F2_1_1  , Final_51_F2_1_1  );
OneRegister RAM_OUT_51_F2_1_2   ( clk , write2_51  , RELUout_F2_1_2  , Final_51_F2_1_2  );
OneRegister RAM_OUT_51_F2_2_1   ( clk , write2_51  , RELUout_F2_2_1  , Final_51_F2_2_1  );
OneRegister RAM_OUT_51_F2_2_2   ( clk , write2_51  , RELUout_F2_2_2  , Final_51_F2_2_2  );
OneRegister RAM_OUT_51_F3_1_1   ( clk , write2_51  , RELUout_F3_1_1  , Final_51_F3_1_1  );
OneRegister RAM_OUT_51_F3_1_2   ( clk , write2_51  , RELUout_F3_1_2  , Final_51_F3_1_2  );
OneRegister RAM_OUT_51_F3_2_1   ( clk , write2_51  , RELUout_F3_2_1  , Final_51_F3_2_1  );
OneRegister RAM_OUT_51_F3_2_2   ( clk , write2_51  , RELUout_F3_2_2  , Final_51_F3_2_2  );
OneRegister RAM_OUT_51_F4_1_1   ( clk , write2_51  , RELUout_F4_1_1  , Final_51_F4_1_1  );
OneRegister RAM_OUT_51_F4_1_2   ( clk , write2_51  , RELUout_F4_1_2  , Final_51_F4_1_2  );
OneRegister RAM_OUT_51_F4_2_1   ( clk , write2_51  , RELUout_F4_2_1  , Final_51_F4_2_1  );
OneRegister RAM_OUT_51_F4_2_2   ( clk , write2_51  , RELUout_F4_2_2  , Final_51_F4_2_2  );
OneRegister RAM_OUT_52_F1_1_1   ( clk , write2_52  , RELUout_F1_1_1  , Final_52_F1_1_1  );
OneRegister RAM_OUT_52_F1_1_2   ( clk , write2_52  , RELUout_F1_1_2  , Final_52_F1_1_2  );
OneRegister RAM_OUT_52_F1_2_1   ( clk , write2_52  , RELUout_F1_2_1  , Final_52_F1_2_1  );
OneRegister RAM_OUT_52_F1_2_2   ( clk , write2_52  , RELUout_F1_2_2  , Final_52_F1_2_2  );
OneRegister RAM_OUT_52_F2_1_1   ( clk , write2_52  , RELUout_F2_1_1  , Final_52_F2_1_1  );
OneRegister RAM_OUT_52_F2_1_2   ( clk , write2_52  , RELUout_F2_1_2  , Final_52_F2_1_2  );
OneRegister RAM_OUT_52_F2_2_1   ( clk , write2_52  , RELUout_F2_2_1  , Final_52_F2_2_1  );
OneRegister RAM_OUT_52_F2_2_2   ( clk , write2_52  , RELUout_F2_2_2  , Final_52_F2_2_2  );
OneRegister RAM_OUT_52_F3_1_1   ( clk , write2_52  , RELUout_F3_1_1  , Final_52_F3_1_1  );
OneRegister RAM_OUT_52_F3_1_2   ( clk , write2_52  , RELUout_F3_1_2  , Final_52_F3_1_2  );
OneRegister RAM_OUT_52_F3_2_1   ( clk , write2_52  , RELUout_F3_2_1  , Final_52_F3_2_1  );
OneRegister RAM_OUT_52_F3_2_2   ( clk , write2_52  , RELUout_F3_2_2  , Final_52_F3_2_2  );
OneRegister RAM_OUT_52_F4_1_1   ( clk , write2_52  , RELUout_F4_1_1  , Final_52_F4_1_1  );
OneRegister RAM_OUT_52_F4_1_2   ( clk , write2_52  , RELUout_F4_1_2  , Final_52_F4_1_2  );
OneRegister RAM_OUT_52_F4_2_1   ( clk , write2_52  , RELUout_F4_2_1  , Final_52_F4_2_1  );
OneRegister RAM_OUT_52_F4_2_2   ( clk , write2_52  , RELUout_F4_2_2  , Final_52_F4_2_2  );
OneRegister RAM_OUT_53_F1_1_1   ( clk , write2_53  , RELUout_F1_1_1  , Final_53_F1_1_1  );
OneRegister RAM_OUT_53_F1_1_2   ( clk , write2_53  , RELUout_F1_1_2  , Final_53_F1_1_2  );
OneRegister RAM_OUT_53_F1_2_1   ( clk , write2_53  , RELUout_F1_2_1  , Final_53_F1_2_1  );
OneRegister RAM_OUT_53_F1_2_2   ( clk , write2_53  , RELUout_F1_2_2  , Final_53_F1_2_2  );
OneRegister RAM_OUT_53_F2_1_1   ( clk , write2_53  , RELUout_F2_1_1  , Final_53_F2_1_1  );
OneRegister RAM_OUT_53_F2_1_2   ( clk , write2_53  , RELUout_F2_1_2  , Final_53_F2_1_2  );
OneRegister RAM_OUT_53_F2_2_1   ( clk , write2_53  , RELUout_F2_2_1  , Final_53_F2_2_1  );
OneRegister RAM_OUT_53_F2_2_2   ( clk , write2_53  , RELUout_F2_2_2  , Final_53_F2_2_2  );
OneRegister RAM_OUT_53_F3_1_1   ( clk , write2_53  , RELUout_F3_1_1  , Final_53_F3_1_1  );
OneRegister RAM_OUT_53_F3_1_2   ( clk , write2_53  , RELUout_F3_1_2  , Final_53_F3_1_2  );
OneRegister RAM_OUT_53_F3_2_1   ( clk , write2_53  , RELUout_F3_2_1  , Final_53_F3_2_1  );
OneRegister RAM_OUT_53_F3_2_2   ( clk , write2_53  , RELUout_F3_2_2  , Final_53_F3_2_2  );
OneRegister RAM_OUT_53_F4_1_1   ( clk , write2_53  , RELUout_F4_1_1  , Final_53_F4_1_1  );
OneRegister RAM_OUT_53_F4_1_2   ( clk , write2_53  , RELUout_F4_1_2  , Final_53_F4_1_2  );
OneRegister RAM_OUT_53_F4_2_1   ( clk , write2_53  , RELUout_F4_2_1  , Final_53_F4_2_1  );
OneRegister RAM_OUT_53_F4_2_2   ( clk , write2_53  , RELUout_F4_2_2  , Final_53_F4_2_2  );
OneRegister RAM_OUT_54_F1_1_1   ( clk , write2_54  , RELUout_F1_1_1  , Final_54_F1_1_1  );
OneRegister RAM_OUT_54_F1_1_2   ( clk , write2_54  , RELUout_F1_1_2  , Final_54_F1_1_2  );
OneRegister RAM_OUT_54_F1_2_1   ( clk , write2_54  , RELUout_F1_2_1  , Final_54_F1_2_1  );
OneRegister RAM_OUT_54_F1_2_2   ( clk , write2_54  , RELUout_F1_2_2  , Final_54_F1_2_2  );
OneRegister RAM_OUT_54_F2_1_1   ( clk , write2_54  , RELUout_F2_1_1  , Final_54_F2_1_1  );
OneRegister RAM_OUT_54_F2_1_2   ( clk , write2_54  , RELUout_F2_1_2  , Final_54_F2_1_2  );
OneRegister RAM_OUT_54_F2_2_1   ( clk , write2_54  , RELUout_F2_2_1  , Final_54_F2_2_1  );
OneRegister RAM_OUT_54_F2_2_2   ( clk , write2_54  , RELUout_F2_2_2  , Final_54_F2_2_2  );
OneRegister RAM_OUT_54_F3_1_1   ( clk , write2_54  , RELUout_F3_1_1  , Final_54_F3_1_1  );
OneRegister RAM_OUT_54_F3_1_2   ( clk , write2_54  , RELUout_F3_1_2  , Final_54_F3_1_2  );
OneRegister RAM_OUT_54_F3_2_1   ( clk , write2_54  , RELUout_F3_2_1  , Final_54_F3_2_1  );
OneRegister RAM_OUT_54_F3_2_2   ( clk , write2_54  , RELUout_F3_2_2  , Final_54_F3_2_2  );
OneRegister RAM_OUT_54_F4_1_1   ( clk , write2_54  , RELUout_F4_1_1  , Final_54_F4_1_1  );
OneRegister RAM_OUT_54_F4_1_2   ( clk , write2_54  , RELUout_F4_1_2  , Final_54_F4_1_2  );
OneRegister RAM_OUT_54_F4_2_1   ( clk , write2_54  , RELUout_F4_2_1  , Final_54_F4_2_1  );
OneRegister RAM_OUT_54_F4_2_2   ( clk , write2_54  , RELUout_F4_2_2  , Final_54_F4_2_2  );
OneRegister RAM_OUT_55_F1_1_1   ( clk , write2_55  , RELUout_F1_1_1  , Final_55_F1_1_1  );
OneRegister RAM_OUT_55_F1_1_2   ( clk , write2_55  , RELUout_F1_1_2  , Final_55_F1_1_2  );
OneRegister RAM_OUT_55_F1_2_1   ( clk , write2_55  , RELUout_F1_2_1  , Final_55_F1_2_1  );
OneRegister RAM_OUT_55_F1_2_2   ( clk , write2_55  , RELUout_F1_2_2  , Final_55_F1_2_2  );
OneRegister RAM_OUT_55_F2_1_1   ( clk , write2_55  , RELUout_F2_1_1  , Final_55_F2_1_1  );
OneRegister RAM_OUT_55_F2_1_2   ( clk , write2_55  , RELUout_F2_1_2  , Final_55_F2_1_2  );
OneRegister RAM_OUT_55_F2_2_1   ( clk , write2_55  , RELUout_F2_2_1  , Final_55_F2_2_1  );
OneRegister RAM_OUT_55_F2_2_2   ( clk , write2_55  , RELUout_F2_2_2  , Final_55_F2_2_2  );
OneRegister RAM_OUT_55_F3_1_1   ( clk , write2_55  , RELUout_F3_1_1  , Final_55_F3_1_1  );
OneRegister RAM_OUT_55_F3_1_2   ( clk , write2_55  , RELUout_F3_1_2  , Final_55_F3_1_2  );
OneRegister RAM_OUT_55_F3_2_1   ( clk , write2_55  , RELUout_F3_2_1  , Final_55_F3_2_1  );
OneRegister RAM_OUT_55_F3_2_2   ( clk , write2_55  , RELUout_F3_2_2  , Final_55_F3_2_2  );
OneRegister RAM_OUT_55_F4_1_1   ( clk , write2_55  , RELUout_F4_1_1  , Final_55_F4_1_1  );
OneRegister RAM_OUT_55_F4_1_2   ( clk , write2_55  , RELUout_F4_1_2  , Final_55_F4_1_2  );
OneRegister RAM_OUT_55_F4_2_1   ( clk , write2_55  , RELUout_F4_2_1  , Final_55_F4_2_1  );
OneRegister RAM_OUT_55_F4_2_2   ( clk , write2_55  , RELUout_F4_2_2  , Final_55_F4_2_2  );
OneRegister RAM_OUT_56_F1_1_1   ( clk , write2_56  , RELUout_F1_1_1  , Final_56_F1_1_1  );
OneRegister RAM_OUT_56_F1_1_2   ( clk , write2_56  , RELUout_F1_1_2  , Final_56_F1_1_2  );
OneRegister RAM_OUT_56_F1_2_1   ( clk , write2_56  , RELUout_F1_2_1  , Final_56_F1_2_1  );
OneRegister RAM_OUT_56_F1_2_2   ( clk , write2_56  , RELUout_F1_2_2  , Final_56_F1_2_2  );
OneRegister RAM_OUT_56_F2_1_1   ( clk , write2_56  , RELUout_F2_1_1  , Final_56_F2_1_1  );
OneRegister RAM_OUT_56_F2_1_2   ( clk , write2_56  , RELUout_F2_1_2  , Final_56_F2_1_2  );
OneRegister RAM_OUT_56_F2_2_1   ( clk , write2_56  , RELUout_F2_2_1  , Final_56_F2_2_1  );
OneRegister RAM_OUT_56_F2_2_2   ( clk , write2_56  , RELUout_F2_2_2  , Final_56_F2_2_2  );
OneRegister RAM_OUT_56_F3_1_1   ( clk , write2_56  , RELUout_F3_1_1  , Final_56_F3_1_1  );
OneRegister RAM_OUT_56_F3_1_2   ( clk , write2_56  , RELUout_F3_1_2  , Final_56_F3_1_2  );
OneRegister RAM_OUT_56_F3_2_1   ( clk , write2_56  , RELUout_F3_2_1  , Final_56_F3_2_1  );
OneRegister RAM_OUT_56_F3_2_2   ( clk , write2_56  , RELUout_F3_2_2  , Final_56_F3_2_2  );
OneRegister RAM_OUT_56_F4_1_1   ( clk , write2_56  , RELUout_F4_1_1  , Final_56_F4_1_1  );
OneRegister RAM_OUT_56_F4_1_2   ( clk , write2_56  , RELUout_F4_1_2  , Final_56_F4_1_2  );
OneRegister RAM_OUT_56_F4_2_1   ( clk , write2_56  , RELUout_F4_2_1  , Final_56_F4_2_1  );
OneRegister RAM_OUT_56_F4_2_2   ( clk , write2_56  , RELUout_F4_2_2  , Final_56_F4_2_2  );
OneRegister RAM_OUT_57_F1_1_1   ( clk , write2_57  , RELUout_F1_1_1  , Final_57_F1_1_1  );
OneRegister RAM_OUT_57_F1_1_2   ( clk , write2_57  , RELUout_F1_1_2  , Final_57_F1_1_2  );
OneRegister RAM_OUT_57_F1_2_1   ( clk , write2_57  , RELUout_F1_2_1  , Final_57_F1_2_1  );
OneRegister RAM_OUT_57_F1_2_2   ( clk , write2_57  , RELUout_F1_2_2  , Final_57_F1_2_2  );
OneRegister RAM_OUT_57_F2_1_1   ( clk , write2_57  , RELUout_F2_1_1  , Final_57_F2_1_1  );
OneRegister RAM_OUT_57_F2_1_2   ( clk , write2_57  , RELUout_F2_1_2  , Final_57_F2_1_2  );
OneRegister RAM_OUT_57_F2_2_1   ( clk , write2_57  , RELUout_F2_2_1  , Final_57_F2_2_1  );
OneRegister RAM_OUT_57_F2_2_2   ( clk , write2_57  , RELUout_F2_2_2  , Final_57_F2_2_2  );
OneRegister RAM_OUT_57_F3_1_1   ( clk , write2_57  , RELUout_F3_1_1  , Final_57_F3_1_1  );
OneRegister RAM_OUT_57_F3_1_2   ( clk , write2_57  , RELUout_F3_1_2  , Final_57_F3_1_2  );
OneRegister RAM_OUT_57_F3_2_1   ( clk , write2_57  , RELUout_F3_2_1  , Final_57_F3_2_1  );
OneRegister RAM_OUT_57_F3_2_2   ( clk , write2_57  , RELUout_F3_2_2  , Final_57_F3_2_2  );
OneRegister RAM_OUT_57_F4_1_1   ( clk , write2_57  , RELUout_F4_1_1  , Final_57_F4_1_1  );
OneRegister RAM_OUT_57_F4_1_2   ( clk , write2_57  , RELUout_F4_1_2  , Final_57_F4_1_2  );
OneRegister RAM_OUT_57_F4_2_1   ( clk , write2_57  , RELUout_F4_2_1  , Final_57_F4_2_1  );
OneRegister RAM_OUT_57_F4_2_2   ( clk , write2_57  , RELUout_F4_2_2  , Final_57_F4_2_2  );
OneRegister RAM_OUT_58_F1_1_1   ( clk , write2_58  , RELUout_F1_1_1  , Final_58_F1_1_1  );
OneRegister RAM_OUT_58_F1_1_2   ( clk , write2_58  , RELUout_F1_1_2  , Final_58_F1_1_2  );
OneRegister RAM_OUT_58_F1_2_1   ( clk , write2_58  , RELUout_F1_2_1  , Final_58_F1_2_1  );
OneRegister RAM_OUT_58_F1_2_2   ( clk , write2_58  , RELUout_F1_2_2  , Final_58_F1_2_2  );
OneRegister RAM_OUT_58_F2_1_1   ( clk , write2_58  , RELUout_F2_1_1  , Final_58_F2_1_1  );
OneRegister RAM_OUT_58_F2_1_2   ( clk , write2_58  , RELUout_F2_1_2  , Final_58_F2_1_2  );
OneRegister RAM_OUT_58_F2_2_1   ( clk , write2_58  , RELUout_F2_2_1  , Final_58_F2_2_1  );
OneRegister RAM_OUT_58_F2_2_2   ( clk , write2_58  , RELUout_F2_2_2  , Final_58_F2_2_2  );
OneRegister RAM_OUT_58_F3_1_1   ( clk , write2_58  , RELUout_F3_1_1  , Final_58_F3_1_1  );
OneRegister RAM_OUT_58_F3_1_2   ( clk , write2_58  , RELUout_F3_1_2  , Final_58_F3_1_2  );
OneRegister RAM_OUT_58_F3_2_1   ( clk , write2_58  , RELUout_F3_2_1  , Final_58_F3_2_1  );
OneRegister RAM_OUT_58_F3_2_2   ( clk , write2_58  , RELUout_F3_2_2  , Final_58_F3_2_2  );
OneRegister RAM_OUT_58_F4_1_1   ( clk , write2_58  , RELUout_F4_1_1  , Final_58_F4_1_1  );
OneRegister RAM_OUT_58_F4_1_2   ( clk , write2_58  , RELUout_F4_1_2  , Final_58_F4_1_2  );
OneRegister RAM_OUT_58_F4_2_1   ( clk , write2_58  , RELUout_F4_2_1  , Final_58_F4_2_1  );
OneRegister RAM_OUT_58_F4_2_2   ( clk , write2_58  , RELUout_F4_2_2  , Final_58_F4_2_2  );
OneRegister RAM_OUT_59_F1_1_1   ( clk , write2_59  , RELUout_F1_1_1  , Final_59_F1_1_1  );
OneRegister RAM_OUT_59_F1_1_2   ( clk , write2_59  , RELUout_F1_1_2  , Final_59_F1_1_2  );
OneRegister RAM_OUT_59_F1_2_1   ( clk , write2_59  , RELUout_F1_2_1  , Final_59_F1_2_1  );
OneRegister RAM_OUT_59_F1_2_2   ( clk , write2_59  , RELUout_F1_2_2  , Final_59_F1_2_2  );
OneRegister RAM_OUT_59_F2_1_1   ( clk , write2_59  , RELUout_F2_1_1  , Final_59_F2_1_1  );
OneRegister RAM_OUT_59_F2_1_2   ( clk , write2_59  , RELUout_F2_1_2  , Final_59_F2_1_2  );
OneRegister RAM_OUT_59_F2_2_1   ( clk , write2_59  , RELUout_F2_2_1  , Final_59_F2_2_1  );
OneRegister RAM_OUT_59_F2_2_2   ( clk , write2_59  , RELUout_F2_2_2  , Final_59_F2_2_2  );
OneRegister RAM_OUT_59_F3_1_1   ( clk , write2_59  , RELUout_F3_1_1  , Final_59_F3_1_1  );
OneRegister RAM_OUT_59_F3_1_2   ( clk , write2_59  , RELUout_F3_1_2  , Final_59_F3_1_2  );
OneRegister RAM_OUT_59_F3_2_1   ( clk , write2_59  , RELUout_F3_2_1  , Final_59_F3_2_1  );
OneRegister RAM_OUT_59_F3_2_2   ( clk , write2_59  , RELUout_F3_2_2  , Final_59_F3_2_2  );
OneRegister RAM_OUT_59_F4_1_1   ( clk , write2_59  , RELUout_F4_1_1  , Final_59_F4_1_1  );
OneRegister RAM_OUT_59_F4_1_2   ( clk , write2_59  , RELUout_F4_1_2  , Final_59_F4_1_2  );
OneRegister RAM_OUT_59_F4_2_1   ( clk , write2_59  , RELUout_F4_2_1  , Final_59_F4_2_1  );
OneRegister RAM_OUT_59_F4_2_2   ( clk , write2_59  , RELUout_F4_2_2  , Final_59_F4_2_2  );
OneRegister RAM_OUT_60_F1_1_1   ( clk , write2_60  , RELUout_F1_1_1  , Final_60_F1_1_1  );
OneRegister RAM_OUT_60_F1_1_2   ( clk , write2_60  , RELUout_F1_1_2  , Final_60_F1_1_2  );
OneRegister RAM_OUT_60_F1_2_1   ( clk , write2_60  , RELUout_F1_2_1  , Final_60_F1_2_1  );
OneRegister RAM_OUT_60_F1_2_2   ( clk , write2_60  , RELUout_F1_2_2  , Final_60_F1_2_2  );
OneRegister RAM_OUT_60_F2_1_1   ( clk , write2_60  , RELUout_F2_1_1  , Final_60_F2_1_1  );
OneRegister RAM_OUT_60_F2_1_2   ( clk , write2_60  , RELUout_F2_1_2  , Final_60_F2_1_2  );
OneRegister RAM_OUT_60_F2_2_1   ( clk , write2_60  , RELUout_F2_2_1  , Final_60_F2_2_1  );
OneRegister RAM_OUT_60_F2_2_2   ( clk , write2_60  , RELUout_F2_2_2  , Final_60_F2_2_2  );
OneRegister RAM_OUT_60_F3_1_1   ( clk , write2_60  , RELUout_F3_1_1  , Final_60_F3_1_1  );
OneRegister RAM_OUT_60_F3_1_2   ( clk , write2_60  , RELUout_F3_1_2  , Final_60_F3_1_2  );
OneRegister RAM_OUT_60_F3_2_1   ( clk , write2_60  , RELUout_F3_2_1  , Final_60_F3_2_1  );
OneRegister RAM_OUT_60_F3_2_2   ( clk , write2_60  , RELUout_F3_2_2  , Final_60_F3_2_2  );
OneRegister RAM_OUT_60_F4_1_1   ( clk , write2_60  , RELUout_F4_1_1  , Final_60_F4_1_1  );
OneRegister RAM_OUT_60_F4_1_2   ( clk , write2_60  , RELUout_F4_1_2  , Final_60_F4_1_2  );
OneRegister RAM_OUT_60_F4_2_1   ( clk , write2_60  , RELUout_F4_2_1  , Final_60_F4_2_1  );
OneRegister RAM_OUT_60_F4_2_2   ( clk , write2_60  , RELUout_F4_2_2  , Final_60_F4_2_2  );
OneRegister RAM_OUT_61_F1_1_1   ( clk , write2_61  , RELUout_F1_1_1  , Final_61_F1_1_1  );
OneRegister RAM_OUT_61_F1_1_2   ( clk , write2_61  , RELUout_F1_1_2  , Final_61_F1_1_2  );
OneRegister RAM_OUT_61_F1_2_1   ( clk , write2_61  , RELUout_F1_2_1  , Final_61_F1_2_1  );
OneRegister RAM_OUT_61_F1_2_2   ( clk , write2_61  , RELUout_F1_2_2  , Final_61_F1_2_2  );
OneRegister RAM_OUT_61_F2_1_1   ( clk , write2_61  , RELUout_F2_1_1  , Final_61_F2_1_1  );
OneRegister RAM_OUT_61_F2_1_2   ( clk , write2_61  , RELUout_F2_1_2  , Final_61_F2_1_2  );
OneRegister RAM_OUT_61_F2_2_1   ( clk , write2_61  , RELUout_F2_2_1  , Final_61_F2_2_1  );
OneRegister RAM_OUT_61_F2_2_2   ( clk , write2_61  , RELUout_F2_2_2  , Final_61_F2_2_2  );
OneRegister RAM_OUT_61_F3_1_1   ( clk , write2_61  , RELUout_F3_1_1  , Final_61_F3_1_1  );
OneRegister RAM_OUT_61_F3_1_2   ( clk , write2_61  , RELUout_F3_1_2  , Final_61_F3_1_2  );
OneRegister RAM_OUT_61_F3_2_1   ( clk , write2_61  , RELUout_F3_2_1  , Final_61_F3_2_1  );
OneRegister RAM_OUT_61_F3_2_2   ( clk , write2_61  , RELUout_F3_2_2  , Final_61_F3_2_2  );
OneRegister RAM_OUT_61_F4_1_1   ( clk , write2_61  , RELUout_F4_1_1  , Final_61_F4_1_1  );
OneRegister RAM_OUT_61_F4_1_2   ( clk , write2_61  , RELUout_F4_1_2  , Final_61_F4_1_2  );
OneRegister RAM_OUT_61_F4_2_1   ( clk , write2_61  , RELUout_F4_2_1  , Final_61_F4_2_1  );
OneRegister RAM_OUT_61_F4_2_2   ( clk , write2_61  , RELUout_F4_2_2  , Final_61_F4_2_2  );
OneRegister RAM_OUT_62_F1_1_1   ( clk , write2_62  , RELUout_F1_1_1  , Final_62_F1_1_1  );
OneRegister RAM_OUT_62_F1_1_2   ( clk , write2_62  , RELUout_F1_1_2  , Final_62_F1_1_2  );
OneRegister RAM_OUT_62_F1_2_1   ( clk , write2_62  , RELUout_F1_2_1  , Final_62_F1_2_1  );
OneRegister RAM_OUT_62_F1_2_2   ( clk , write2_62  , RELUout_F1_2_2  , Final_62_F1_2_2  );
OneRegister RAM_OUT_62_F2_1_1   ( clk , write2_62  , RELUout_F2_1_1  , Final_62_F2_1_1  );
OneRegister RAM_OUT_62_F2_1_2   ( clk , write2_62  , RELUout_F2_1_2  , Final_62_F2_1_2  );
OneRegister RAM_OUT_62_F2_2_1   ( clk , write2_62  , RELUout_F2_2_1  , Final_62_F2_2_1  );
OneRegister RAM_OUT_62_F2_2_2   ( clk , write2_62  , RELUout_F2_2_2  , Final_62_F2_2_2  );
OneRegister RAM_OUT_62_F3_1_1   ( clk , write2_62  , RELUout_F3_1_1  , Final_62_F3_1_1  );
OneRegister RAM_OUT_62_F3_1_2   ( clk , write2_62  , RELUout_F3_1_2  , Final_62_F3_1_2  );
OneRegister RAM_OUT_62_F3_2_1   ( clk , write2_62  , RELUout_F3_2_1  , Final_62_F3_2_1  );
OneRegister RAM_OUT_62_F3_2_2   ( clk , write2_62  , RELUout_F3_2_2  , Final_62_F3_2_2  );
OneRegister RAM_OUT_62_F4_1_1   ( clk , write2_62  , RELUout_F4_1_1  , Final_62_F4_1_1  );
OneRegister RAM_OUT_62_F4_1_2   ( clk , write2_62  , RELUout_F4_1_2  , Final_62_F4_1_2  );
OneRegister RAM_OUT_62_F4_2_1   ( clk , write2_62  , RELUout_F4_2_1  , Final_62_F4_2_1  );
OneRegister RAM_OUT_62_F4_2_2   ( clk , write2_62  , RELUout_F4_2_2  , Final_62_F4_2_2  );
OneRegister RAM_OUT_63_F1_1_1   ( clk , write2_63  , RELUout_F1_1_1  , Final_63_F1_1_1  );
OneRegister RAM_OUT_63_F1_1_2   ( clk , write2_63  , RELUout_F1_1_2  , Final_63_F1_1_2  );
OneRegister RAM_OUT_63_F1_2_1   ( clk , write2_63  , RELUout_F1_2_1  , Final_63_F1_2_1  );
OneRegister RAM_OUT_63_F1_2_2   ( clk , write2_63  , RELUout_F1_2_2  , Final_63_F1_2_2  );
OneRegister RAM_OUT_63_F2_1_1   ( clk , write2_63  , RELUout_F2_1_1  , Final_63_F2_1_1  );
OneRegister RAM_OUT_63_F2_1_2   ( clk , write2_63  , RELUout_F2_1_2  , Final_63_F2_1_2  );
OneRegister RAM_OUT_63_F2_2_1   ( clk , write2_63  , RELUout_F2_2_1  , Final_63_F2_2_1  );
OneRegister RAM_OUT_63_F2_2_2   ( clk , write2_63  , RELUout_F2_2_2  , Final_63_F2_2_2  );
OneRegister RAM_OUT_63_F3_1_1   ( clk , write2_63  , RELUout_F3_1_1  , Final_63_F3_1_1  );
OneRegister RAM_OUT_63_F3_1_2   ( clk , write2_63  , RELUout_F3_1_2  , Final_63_F3_1_2  );
OneRegister RAM_OUT_63_F3_2_1   ( clk , write2_63  , RELUout_F3_2_1  , Final_63_F3_2_1  );
OneRegister RAM_OUT_63_F3_2_2   ( clk , write2_63  , RELUout_F3_2_2  , Final_63_F3_2_2  );
OneRegister RAM_OUT_63_F4_1_1   ( clk , write2_63  , RELUout_F4_1_1  , Final_63_F4_1_1  );
OneRegister RAM_OUT_63_F4_1_2   ( clk , write2_63  , RELUout_F4_1_2  , Final_63_F4_1_2  );
OneRegister RAM_OUT_63_F4_2_1   ( clk , write2_63  , RELUout_F4_2_1  , Final_63_F4_2_1  );
OneRegister RAM_OUT_63_F4_2_2   ( clk , write2_63  , RELUout_F4_2_2  , Final_63_F4_2_2  );
OneRegister RAM_OUT_64_F1_1_1   ( clk , write2_64  , RELUout_F1_1_1  , Final_64_F1_1_1  );
OneRegister RAM_OUT_64_F1_1_2   ( clk , write2_64  , RELUout_F1_1_2  , Final_64_F1_1_2  );
OneRegister RAM_OUT_64_F1_2_1   ( clk , write2_64  , RELUout_F1_2_1  , Final_64_F1_2_1  );
OneRegister RAM_OUT_64_F1_2_2   ( clk , write2_64  , RELUout_F1_2_2  , Final_64_F1_2_2  );
OneRegister RAM_OUT_64_F2_1_1   ( clk , write2_64  , RELUout_F2_1_1  , Final_64_F2_1_1  );
OneRegister RAM_OUT_64_F2_1_2   ( clk , write2_64  , RELUout_F2_1_2  , Final_64_F2_1_2  );
OneRegister RAM_OUT_64_F2_2_1   ( clk , write2_64  , RELUout_F2_2_1  , Final_64_F2_2_1  );
OneRegister RAM_OUT_64_F2_2_2   ( clk , write2_64  , RELUout_F2_2_2  , Final_64_F2_2_2  );
OneRegister RAM_OUT_64_F3_1_1   ( clk , write2_64  , RELUout_F3_1_1  , Final_64_F3_1_1  );
OneRegister RAM_OUT_64_F3_1_2   ( clk , write2_64  , RELUout_F3_1_2  , Final_64_F3_1_2  );
OneRegister RAM_OUT_64_F3_2_1   ( clk , write2_64  , RELUout_F3_2_1  , Final_64_F3_2_1  );
OneRegister RAM_OUT_64_F3_2_2   ( clk , write2_64  , RELUout_F3_2_2  , Final_64_F3_2_2  );
OneRegister RAM_OUT_64_F4_1_1   ( clk , write2_64  , RELUout_F4_1_1  , Final_64_F4_1_1  );
OneRegister RAM_OUT_64_F4_1_2   ( clk , write2_64  , RELUout_F4_1_2  , Final_64_F4_1_2  );
OneRegister RAM_OUT_64_F4_2_1   ( clk , write2_64  , RELUout_F4_2_1  , Final_64_F4_2_1  );
OneRegister RAM_OUT_64_F4_2_2   ( clk , write2_64  , RELUout_F4_2_2  , Final_64_F4_2_2  );
OneRegister RAM_OUT_65_F1_1_1   ( clk , write2_65  , RELUout_F1_1_1  , Final_65_F1_1_1  );
OneRegister RAM_OUT_65_F1_1_2   ( clk , write2_65  , RELUout_F1_1_2  , Final_65_F1_1_2  );
OneRegister RAM_OUT_65_F1_2_1   ( clk , write2_65  , RELUout_F1_2_1  , Final_65_F1_2_1  );
OneRegister RAM_OUT_65_F1_2_2   ( clk , write2_65  , RELUout_F1_2_2  , Final_65_F1_2_2  );
OneRegister RAM_OUT_65_F2_1_1   ( clk , write2_65  , RELUout_F2_1_1  , Final_65_F2_1_1  );
OneRegister RAM_OUT_65_F2_1_2   ( clk , write2_65  , RELUout_F2_1_2  , Final_65_F2_1_2  );
OneRegister RAM_OUT_65_F2_2_1   ( clk , write2_65  , RELUout_F2_2_1  , Final_65_F2_2_1  );
OneRegister RAM_OUT_65_F2_2_2   ( clk , write2_65  , RELUout_F2_2_2  , Final_65_F2_2_2  );
OneRegister RAM_OUT_65_F3_1_1   ( clk , write2_65  , RELUout_F3_1_1  , Final_65_F3_1_1  );
OneRegister RAM_OUT_65_F3_1_2   ( clk , write2_65  , RELUout_F3_1_2  , Final_65_F3_1_2  );
OneRegister RAM_OUT_65_F3_2_1   ( clk , write2_65  , RELUout_F3_2_1  , Final_65_F3_2_1  );
OneRegister RAM_OUT_65_F3_2_2   ( clk , write2_65  , RELUout_F3_2_2  , Final_65_F3_2_2  );
OneRegister RAM_OUT_65_F4_1_1   ( clk , write2_65  , RELUout_F4_1_1  , Final_65_F4_1_1  );
OneRegister RAM_OUT_65_F4_1_2   ( clk , write2_65  , RELUout_F4_1_2  , Final_65_F4_1_2  );
OneRegister RAM_OUT_65_F4_2_1   ( clk , write2_65  , RELUout_F4_2_1  , Final_65_F4_2_1  );
OneRegister RAM_OUT_65_F4_2_2   ( clk , write2_65  , RELUout_F4_2_2  , Final_65_F4_2_2  );
OneRegister RAM_OUT_66_F1_1_1   ( clk , write2_66  , RELUout_F1_1_1  , Final_66_F1_1_1  );
OneRegister RAM_OUT_66_F1_1_2   ( clk , write2_66  , RELUout_F1_1_2  , Final_66_F1_1_2  );
OneRegister RAM_OUT_66_F1_2_1   ( clk , write2_66  , RELUout_F1_2_1  , Final_66_F1_2_1  );
OneRegister RAM_OUT_66_F1_2_2   ( clk , write2_66  , RELUout_F1_2_2  , Final_66_F1_2_2  );
OneRegister RAM_OUT_66_F2_1_1   ( clk , write2_66  , RELUout_F2_1_1  , Final_66_F2_1_1  );
OneRegister RAM_OUT_66_F2_1_2   ( clk , write2_66  , RELUout_F2_1_2  , Final_66_F2_1_2  );
OneRegister RAM_OUT_66_F2_2_1   ( clk , write2_66  , RELUout_F2_2_1  , Final_66_F2_2_1  );
OneRegister RAM_OUT_66_F2_2_2   ( clk , write2_66  , RELUout_F2_2_2  , Final_66_F2_2_2  );
OneRegister RAM_OUT_66_F3_1_1   ( clk , write2_66  , RELUout_F3_1_1  , Final_66_F3_1_1  );
OneRegister RAM_OUT_66_F3_1_2   ( clk , write2_66  , RELUout_F3_1_2  , Final_66_F3_1_2  );
OneRegister RAM_OUT_66_F3_2_1   ( clk , write2_66  , RELUout_F3_2_1  , Final_66_F3_2_1  );
OneRegister RAM_OUT_66_F3_2_2   ( clk , write2_66  , RELUout_F3_2_2  , Final_66_F3_2_2  );
OneRegister RAM_OUT_66_F4_1_1   ( clk , write2_66  , RELUout_F4_1_1  , Final_66_F4_1_1  );
OneRegister RAM_OUT_66_F4_1_2   ( clk , write2_66  , RELUout_F4_1_2  , Final_66_F4_1_2  );
OneRegister RAM_OUT_66_F4_2_1   ( clk , write2_66  , RELUout_F4_2_1  , Final_66_F4_2_1  );
OneRegister RAM_OUT_66_F4_2_2   ( clk , write2_66  , RELUout_F4_2_2  , Final_66_F4_2_2  );
OneRegister RAM_OUT_67_F1_1_1   ( clk , write2_67  , RELUout_F1_1_1  , Final_67_F1_1_1  );
OneRegister RAM_OUT_67_F1_1_2   ( clk , write2_67  , RELUout_F1_1_2  , Final_67_F1_1_2  );
OneRegister RAM_OUT_67_F1_2_1   ( clk , write2_67  , RELUout_F1_2_1  , Final_67_F1_2_1  );
OneRegister RAM_OUT_67_F1_2_2   ( clk , write2_67  , RELUout_F1_2_2  , Final_67_F1_2_2  );
OneRegister RAM_OUT_67_F2_1_1   ( clk , write2_67  , RELUout_F2_1_1  , Final_67_F2_1_1  );
OneRegister RAM_OUT_67_F2_1_2   ( clk , write2_67  , RELUout_F2_1_2  , Final_67_F2_1_2  );
OneRegister RAM_OUT_67_F2_2_1   ( clk , write2_67  , RELUout_F2_2_1  , Final_67_F2_2_1  );
OneRegister RAM_OUT_67_F2_2_2   ( clk , write2_67  , RELUout_F2_2_2  , Final_67_F2_2_2  );
OneRegister RAM_OUT_67_F3_1_1   ( clk , write2_67  , RELUout_F3_1_1  , Final_67_F3_1_1  );
OneRegister RAM_OUT_67_F3_1_2   ( clk , write2_67  , RELUout_F3_1_2  , Final_67_F3_1_2  );
OneRegister RAM_OUT_67_F3_2_1   ( clk , write2_67  , RELUout_F3_2_1  , Final_67_F3_2_1  );
OneRegister RAM_OUT_67_F3_2_2   ( clk , write2_67  , RELUout_F3_2_2  , Final_67_F3_2_2  );
OneRegister RAM_OUT_67_F4_1_1   ( clk , write2_67  , RELUout_F4_1_1  , Final_67_F4_1_1  );
OneRegister RAM_OUT_67_F4_1_2   ( clk , write2_67  , RELUout_F4_1_2  , Final_67_F4_1_2  );
OneRegister RAM_OUT_67_F4_2_1   ( clk , write2_67  , RELUout_F4_2_1  , Final_67_F4_2_1  );
OneRegister RAM_OUT_67_F4_2_2   ( clk , write2_67  , RELUout_F4_2_2  , Final_67_F4_2_2  );
OneRegister RAM_OUT_68_F1_1_1   ( clk , write2_68  , RELUout_F1_1_1  , Final_68_F1_1_1  );
OneRegister RAM_OUT_68_F1_1_2   ( clk , write2_68  , RELUout_F1_1_2  , Final_68_F1_1_2  );
OneRegister RAM_OUT_68_F1_2_1   ( clk , write2_68  , RELUout_F1_2_1  , Final_68_F1_2_1  );
OneRegister RAM_OUT_68_F1_2_2   ( clk , write2_68  , RELUout_F1_2_2  , Final_68_F1_2_2  );
OneRegister RAM_OUT_68_F2_1_1   ( clk , write2_68  , RELUout_F2_1_1  , Final_68_F2_1_1  );
OneRegister RAM_OUT_68_F2_1_2   ( clk , write2_68  , RELUout_F2_1_2  , Final_68_F2_1_2  );
OneRegister RAM_OUT_68_F2_2_1   ( clk , write2_68  , RELUout_F2_2_1  , Final_68_F2_2_1  );
OneRegister RAM_OUT_68_F2_2_2   ( clk , write2_68  , RELUout_F2_2_2  , Final_68_F2_2_2  );
OneRegister RAM_OUT_68_F3_1_1   ( clk , write2_68  , RELUout_F3_1_1  , Final_68_F3_1_1  );
OneRegister RAM_OUT_68_F3_1_2   ( clk , write2_68  , RELUout_F3_1_2  , Final_68_F3_1_2  );
OneRegister RAM_OUT_68_F3_2_1   ( clk , write2_68  , RELUout_F3_2_1  , Final_68_F3_2_1  );
OneRegister RAM_OUT_68_F3_2_2   ( clk , write2_68  , RELUout_F3_2_2  , Final_68_F3_2_2  );
OneRegister RAM_OUT_68_F4_1_1   ( clk , write2_68  , RELUout_F4_1_1  , Final_68_F4_1_1  );
OneRegister RAM_OUT_68_F4_1_2   ( clk , write2_68  , RELUout_F4_1_2  , Final_68_F4_1_2  );
OneRegister RAM_OUT_68_F4_2_1   ( clk , write2_68  , RELUout_F4_2_1  , Final_68_F4_2_1  );
OneRegister RAM_OUT_68_F4_2_2   ( clk , write2_68  , RELUout_F4_2_2  , Final_68_F4_2_2  );
OneRegister RAM_OUT_69_F1_1_1   ( clk , write2_69  , RELUout_F1_1_1  , Final_69_F1_1_1  );
OneRegister RAM_OUT_69_F1_1_2   ( clk , write2_69  , RELUout_F1_1_2  , Final_69_F1_1_2  );
OneRegister RAM_OUT_69_F1_2_1   ( clk , write2_69  , RELUout_F1_2_1  , Final_69_F1_2_1  );
OneRegister RAM_OUT_69_F1_2_2   ( clk , write2_69  , RELUout_F1_2_2  , Final_69_F1_2_2  );
OneRegister RAM_OUT_69_F2_1_1   ( clk , write2_69  , RELUout_F2_1_1  , Final_69_F2_1_1  );
OneRegister RAM_OUT_69_F2_1_2   ( clk , write2_69  , RELUout_F2_1_2  , Final_69_F2_1_2  );
OneRegister RAM_OUT_69_F2_2_1   ( clk , write2_69  , RELUout_F2_2_1  , Final_69_F2_2_1  );
OneRegister RAM_OUT_69_F2_2_2   ( clk , write2_69  , RELUout_F2_2_2  , Final_69_F2_2_2  );
OneRegister RAM_OUT_69_F3_1_1   ( clk , write2_69  , RELUout_F3_1_1  , Final_69_F3_1_1  );
OneRegister RAM_OUT_69_F3_1_2   ( clk , write2_69  , RELUout_F3_1_2  , Final_69_F3_1_2  );
OneRegister RAM_OUT_69_F3_2_1   ( clk , write2_69  , RELUout_F3_2_1  , Final_69_F3_2_1  );
OneRegister RAM_OUT_69_F3_2_2   ( clk , write2_69  , RELUout_F3_2_2  , Final_69_F3_2_2  );
OneRegister RAM_OUT_69_F4_1_1   ( clk , write2_69  , RELUout_F4_1_1  , Final_69_F4_1_1  );
OneRegister RAM_OUT_69_F4_1_2   ( clk , write2_69  , RELUout_F4_1_2  , Final_69_F4_1_2  );
OneRegister RAM_OUT_69_F4_2_1   ( clk , write2_69  , RELUout_F4_2_1  , Final_69_F4_2_1  );
OneRegister RAM_OUT_69_F4_2_2   ( clk , write2_69  , RELUout_F4_2_2  , Final_69_F4_2_2  );
OneRegister RAM_OUT_70_F1_1_1   ( clk , write2_70  , RELUout_F1_1_1  , Final_70_F1_1_1  );
OneRegister RAM_OUT_70_F1_1_2   ( clk , write2_70  , RELUout_F1_1_2  , Final_70_F1_1_2  );
OneRegister RAM_OUT_70_F1_2_1   ( clk , write2_70  , RELUout_F1_2_1  , Final_70_F1_2_1  );
OneRegister RAM_OUT_70_F1_2_2   ( clk , write2_70  , RELUout_F1_2_2  , Final_70_F1_2_2  );
OneRegister RAM_OUT_70_F2_1_1   ( clk , write2_70  , RELUout_F2_1_1  , Final_70_F2_1_1  );
OneRegister RAM_OUT_70_F2_1_2   ( clk , write2_70  , RELUout_F2_1_2  , Final_70_F2_1_2  );
OneRegister RAM_OUT_70_F2_2_1   ( clk , write2_70  , RELUout_F2_2_1  , Final_70_F2_2_1  );
OneRegister RAM_OUT_70_F2_2_2   ( clk , write2_70  , RELUout_F2_2_2  , Final_70_F2_2_2  );
OneRegister RAM_OUT_70_F3_1_1   ( clk , write2_70  , RELUout_F3_1_1  , Final_70_F3_1_1  );
OneRegister RAM_OUT_70_F3_1_2   ( clk , write2_70  , RELUout_F3_1_2  , Final_70_F3_1_2  );
OneRegister RAM_OUT_70_F3_2_1   ( clk , write2_70  , RELUout_F3_2_1  , Final_70_F3_2_1  );
OneRegister RAM_OUT_70_F3_2_2   ( clk , write2_70  , RELUout_F3_2_2  , Final_70_F3_2_2  );
OneRegister RAM_OUT_70_F4_1_1   ( clk , write2_70  , RELUout_F4_1_1  , Final_70_F4_1_1  );
OneRegister RAM_OUT_70_F4_1_2   ( clk , write2_70  , RELUout_F4_1_2  , Final_70_F4_1_2  );
OneRegister RAM_OUT_70_F4_2_1   ( clk , write2_70  , RELUout_F4_2_1  , Final_70_F4_2_1  );
OneRegister RAM_OUT_70_F4_2_2   ( clk , write2_70  , RELUout_F4_2_2  , Final_70_F4_2_2  );
OneRegister RAM_OUT_71_F1_1_1   ( clk , write2_71  , RELUout_F1_1_1  , Final_71_F1_1_1  );
OneRegister RAM_OUT_71_F1_1_2   ( clk , write2_71  , RELUout_F1_1_2  , Final_71_F1_1_2  );
OneRegister RAM_OUT_71_F1_2_1   ( clk , write2_71  , RELUout_F1_2_1  , Final_71_F1_2_1  );
OneRegister RAM_OUT_71_F1_2_2   ( clk , write2_71  , RELUout_F1_2_2  , Final_71_F1_2_2  );
OneRegister RAM_OUT_71_F2_1_1   ( clk , write2_71  , RELUout_F2_1_1  , Final_71_F2_1_1  );
OneRegister RAM_OUT_71_F2_1_2   ( clk , write2_71  , RELUout_F2_1_2  , Final_71_F2_1_2  );
OneRegister RAM_OUT_71_F2_2_1   ( clk , write2_71  , RELUout_F2_2_1  , Final_71_F2_2_1  );
OneRegister RAM_OUT_71_F2_2_2   ( clk , write2_71  , RELUout_F2_2_2  , Final_71_F2_2_2  );
OneRegister RAM_OUT_71_F3_1_1   ( clk , write2_71  , RELUout_F3_1_1  , Final_71_F3_1_1  );
OneRegister RAM_OUT_71_F3_1_2   ( clk , write2_71  , RELUout_F3_1_2  , Final_71_F3_1_2  );
OneRegister RAM_OUT_71_F3_2_1   ( clk , write2_71  , RELUout_F3_2_1  , Final_71_F3_2_1  );
OneRegister RAM_OUT_71_F3_2_2   ( clk , write2_71  , RELUout_F3_2_2  , Final_71_F3_2_2  );
OneRegister RAM_OUT_71_F4_1_1   ( clk , write2_71  , RELUout_F4_1_1  , Final_71_F4_1_1  );
OneRegister RAM_OUT_71_F4_1_2   ( clk , write2_71  , RELUout_F4_1_2  , Final_71_F4_1_2  );
OneRegister RAM_OUT_71_F4_2_1   ( clk , write2_71  , RELUout_F4_2_1  , Final_71_F4_2_1  );
OneRegister RAM_OUT_71_F4_2_2   ( clk , write2_71  , RELUout_F4_2_2  , Final_71_F4_2_2  );
OneRegister RAM_OUT_72_F1_1_1   ( clk , write2_72  , RELUout_F1_1_1  , Final_72_F1_1_1  );
OneRegister RAM_OUT_72_F1_1_2   ( clk , write2_72  , RELUout_F1_1_2  , Final_72_F1_1_2  );
OneRegister RAM_OUT_72_F1_2_1   ( clk , write2_72  , RELUout_F1_2_1  , Final_72_F1_2_1  );
OneRegister RAM_OUT_72_F1_2_2   ( clk , write2_72  , RELUout_F1_2_2  , Final_72_F1_2_2  );
OneRegister RAM_OUT_72_F2_1_1   ( clk , write2_72  , RELUout_F2_1_1  , Final_72_F2_1_1  );
OneRegister RAM_OUT_72_F2_1_2   ( clk , write2_72  , RELUout_F2_1_2  , Final_72_F2_1_2  );
OneRegister RAM_OUT_72_F2_2_1   ( clk , write2_72  , RELUout_F2_2_1  , Final_72_F2_2_1  );
OneRegister RAM_OUT_72_F2_2_2   ( clk , write2_72  , RELUout_F2_2_2  , Final_72_F2_2_2  );
OneRegister RAM_OUT_72_F3_1_1   ( clk , write2_72  , RELUout_F3_1_1  , Final_72_F3_1_1  );
OneRegister RAM_OUT_72_F3_1_2   ( clk , write2_72  , RELUout_F3_1_2  , Final_72_F3_1_2  );
OneRegister RAM_OUT_72_F3_2_1   ( clk , write2_72  , RELUout_F3_2_1  , Final_72_F3_2_1  );
OneRegister RAM_OUT_72_F3_2_2   ( clk , write2_72  , RELUout_F3_2_2  , Final_72_F3_2_2  );
OneRegister RAM_OUT_72_F4_1_1   ( clk , write2_72  , RELUout_F4_1_1  , Final_72_F4_1_1  );
OneRegister RAM_OUT_72_F4_1_2   ( clk , write2_72  , RELUout_F4_1_2  , Final_72_F4_1_2  );
OneRegister RAM_OUT_72_F4_2_1   ( clk , write2_72  , RELUout_F4_2_1  , Final_72_F4_2_1  );
OneRegister RAM_OUT_72_F4_2_2   ( clk , write2_72  , RELUout_F4_2_2  , Final_72_F4_2_2  );
OneRegister RAM_OUT_73_F1_1_1   ( clk , write2_73  , RELUout_F1_1_1  , Final_73_F1_1_1  );
OneRegister RAM_OUT_73_F1_1_2   ( clk , write2_73  , RELUout_F1_1_2  , Final_73_F1_1_2  );
OneRegister RAM_OUT_73_F1_2_1   ( clk , write2_73  , RELUout_F1_2_1  , Final_73_F1_2_1  );
OneRegister RAM_OUT_73_F1_2_2   ( clk , write2_73  , RELUout_F1_2_2  , Final_73_F1_2_2  );
OneRegister RAM_OUT_73_F2_1_1   ( clk , write2_73  , RELUout_F2_1_1  , Final_73_F2_1_1  );
OneRegister RAM_OUT_73_F2_1_2   ( clk , write2_73  , RELUout_F2_1_2  , Final_73_F2_1_2  );
OneRegister RAM_OUT_73_F2_2_1   ( clk , write2_73  , RELUout_F2_2_1  , Final_73_F2_2_1  );
OneRegister RAM_OUT_73_F2_2_2   ( clk , write2_73  , RELUout_F2_2_2  , Final_73_F2_2_2  );
OneRegister RAM_OUT_73_F3_1_1   ( clk , write2_73  , RELUout_F3_1_1  , Final_73_F3_1_1  );
OneRegister RAM_OUT_73_F3_1_2   ( clk , write2_73  , RELUout_F3_1_2  , Final_73_F3_1_2  );
OneRegister RAM_OUT_73_F3_2_1   ( clk , write2_73  , RELUout_F3_2_1  , Final_73_F3_2_1  );
OneRegister RAM_OUT_73_F3_2_2   ( clk , write2_73  , RELUout_F3_2_2  , Final_73_F3_2_2  );
OneRegister RAM_OUT_73_F4_1_1   ( clk , write2_73  , RELUout_F4_1_1  , Final_73_F4_1_1  );
OneRegister RAM_OUT_73_F4_1_2   ( clk , write2_73  , RELUout_F4_1_2  , Final_73_F4_1_2  );
OneRegister RAM_OUT_73_F4_2_1   ( clk , write2_73  , RELUout_F4_2_1  , Final_73_F4_2_1  );
OneRegister RAM_OUT_73_F4_2_2   ( clk , write2_73  , RELUout_F4_2_2  , Final_73_F4_2_2  );
OneRegister RAM_OUT_74_F1_1_1   ( clk , write2_74  , RELUout_F1_1_1  , Final_74_F1_1_1  );
OneRegister RAM_OUT_74_F1_1_2   ( clk , write2_74  , RELUout_F1_1_2  , Final_74_F1_1_2  );
OneRegister RAM_OUT_74_F1_2_1   ( clk , write2_74  , RELUout_F1_2_1  , Final_74_F1_2_1  );
OneRegister RAM_OUT_74_F1_2_2   ( clk , write2_74  , RELUout_F1_2_2  , Final_74_F1_2_2  );
OneRegister RAM_OUT_74_F2_1_1   ( clk , write2_74  , RELUout_F2_1_1  , Final_74_F2_1_1  );
OneRegister RAM_OUT_74_F2_1_2   ( clk , write2_74  , RELUout_F2_1_2  , Final_74_F2_1_2  );
OneRegister RAM_OUT_74_F2_2_1   ( clk , write2_74  , RELUout_F2_2_1  , Final_74_F2_2_1  );
OneRegister RAM_OUT_74_F2_2_2   ( clk , write2_74  , RELUout_F2_2_2  , Final_74_F2_2_2  );
OneRegister RAM_OUT_74_F3_1_1   ( clk , write2_74  , RELUout_F3_1_1  , Final_74_F3_1_1  );
OneRegister RAM_OUT_74_F3_1_2   ( clk , write2_74  , RELUout_F3_1_2  , Final_74_F3_1_2  );
OneRegister RAM_OUT_74_F3_2_1   ( clk , write2_74  , RELUout_F3_2_1  , Final_74_F3_2_1  );
OneRegister RAM_OUT_74_F3_2_2   ( clk , write2_74  , RELUout_F3_2_2  , Final_74_F3_2_2  );
OneRegister RAM_OUT_74_F4_1_1   ( clk , write2_74  , RELUout_F4_1_1  , Final_74_F4_1_1  );
OneRegister RAM_OUT_74_F4_1_2   ( clk , write2_74  , RELUout_F4_1_2  , Final_74_F4_1_2  );
OneRegister RAM_OUT_74_F4_2_1   ( clk , write2_74  , RELUout_F4_2_1  , Final_74_F4_2_1  );
OneRegister RAM_OUT_74_F4_2_2   ( clk , write2_74  , RELUout_F4_2_2  , Final_74_F4_2_2  );
OneRegister RAM_OUT_75_F1_1_1   ( clk , write2_75  , RELUout_F1_1_1  , Final_75_F1_1_1  );
OneRegister RAM_OUT_75_F1_1_2   ( clk , write2_75  , RELUout_F1_1_2  , Final_75_F1_1_2  );
OneRegister RAM_OUT_75_F1_2_1   ( clk , write2_75  , RELUout_F1_2_1  , Final_75_F1_2_1  );
OneRegister RAM_OUT_75_F1_2_2   ( clk , write2_75  , RELUout_F1_2_2  , Final_75_F1_2_2  );
OneRegister RAM_OUT_75_F2_1_1   ( clk , write2_75  , RELUout_F2_1_1  , Final_75_F2_1_1  );
OneRegister RAM_OUT_75_F2_1_2   ( clk , write2_75  , RELUout_F2_1_2  , Final_75_F2_1_2  );
OneRegister RAM_OUT_75_F2_2_1   ( clk , write2_75  , RELUout_F2_2_1  , Final_75_F2_2_1  );
OneRegister RAM_OUT_75_F2_2_2   ( clk , write2_75  , RELUout_F2_2_2  , Final_75_F2_2_2  );
OneRegister RAM_OUT_75_F3_1_1   ( clk , write2_75  , RELUout_F3_1_1  , Final_75_F3_1_1  );
OneRegister RAM_OUT_75_F3_1_2   ( clk , write2_75  , RELUout_F3_1_2  , Final_75_F3_1_2  );
OneRegister RAM_OUT_75_F3_2_1   ( clk , write2_75  , RELUout_F3_2_1  , Final_75_F3_2_1  );
OneRegister RAM_OUT_75_F3_2_2   ( clk , write2_75  , RELUout_F3_2_2  , Final_75_F3_2_2  );
OneRegister RAM_OUT_75_F4_1_1   ( clk , write2_75  , RELUout_F4_1_1  , Final_75_F4_1_1  );
OneRegister RAM_OUT_75_F4_1_2   ( clk , write2_75  , RELUout_F4_1_2  , Final_75_F4_1_2  );
OneRegister RAM_OUT_75_F4_2_1   ( clk , write2_75  , RELUout_F4_2_1  , Final_75_F4_2_1  );
OneRegister RAM_OUT_75_F4_2_2   ( clk , write2_75  , RELUout_F4_2_2  , Final_75_F4_2_2  );
OneRegister RAM_OUT_76_F1_1_1   ( clk , write2_76  , RELUout_F1_1_1  , Final_76_F1_1_1  );
OneRegister RAM_OUT_76_F1_1_2   ( clk , write2_76  , RELUout_F1_1_2  , Final_76_F1_1_2  );
OneRegister RAM_OUT_76_F1_2_1   ( clk , write2_76  , RELUout_F1_2_1  , Final_76_F1_2_1  );
OneRegister RAM_OUT_76_F1_2_2   ( clk , write2_76  , RELUout_F1_2_2  , Final_76_F1_2_2  );
OneRegister RAM_OUT_76_F2_1_1   ( clk , write2_76  , RELUout_F2_1_1  , Final_76_F2_1_1  );
OneRegister RAM_OUT_76_F2_1_2   ( clk , write2_76  , RELUout_F2_1_2  , Final_76_F2_1_2  );
OneRegister RAM_OUT_76_F2_2_1   ( clk , write2_76  , RELUout_F2_2_1  , Final_76_F2_2_1  );
OneRegister RAM_OUT_76_F2_2_2   ( clk , write2_76  , RELUout_F2_2_2  , Final_76_F2_2_2  );
OneRegister RAM_OUT_76_F3_1_1   ( clk , write2_76  , RELUout_F3_1_1  , Final_76_F3_1_1  );
OneRegister RAM_OUT_76_F3_1_2   ( clk , write2_76  , RELUout_F3_1_2  , Final_76_F3_1_2  );
OneRegister RAM_OUT_76_F3_2_1   ( clk , write2_76  , RELUout_F3_2_1  , Final_76_F3_2_1  );
OneRegister RAM_OUT_76_F3_2_2   ( clk , write2_76  , RELUout_F3_2_2  , Final_76_F3_2_2  );
OneRegister RAM_OUT_76_F4_1_1   ( clk , write2_76  , RELUout_F4_1_1  , Final_76_F4_1_1  );
OneRegister RAM_OUT_76_F4_1_2   ( clk , write2_76  , RELUout_F4_1_2  , Final_76_F4_1_2  );
OneRegister RAM_OUT_76_F4_2_1   ( clk , write2_76  , RELUout_F4_2_1  , Final_76_F4_2_1  );
OneRegister RAM_OUT_76_F4_2_2   ( clk , write2_76  , RELUout_F4_2_2  , Final_76_F4_2_2  );
OneRegister RAM_OUT_77_F1_1_1   ( clk , write2_77  , RELUout_F1_1_1  , Final_77_F1_1_1  );
OneRegister RAM_OUT_77_F1_1_2   ( clk , write2_77  , RELUout_F1_1_2  , Final_77_F1_1_2  );
OneRegister RAM_OUT_77_F1_2_1   ( clk , write2_77  , RELUout_F1_2_1  , Final_77_F1_2_1  );
OneRegister RAM_OUT_77_F1_2_2   ( clk , write2_77  , RELUout_F1_2_2  , Final_77_F1_2_2  );
OneRegister RAM_OUT_77_F2_1_1   ( clk , write2_77  , RELUout_F2_1_1  , Final_77_F2_1_1  );
OneRegister RAM_OUT_77_F2_1_2   ( clk , write2_77  , RELUout_F2_1_2  , Final_77_F2_1_2  );
OneRegister RAM_OUT_77_F2_2_1   ( clk , write2_77  , RELUout_F2_2_1  , Final_77_F2_2_1  );
OneRegister RAM_OUT_77_F2_2_2   ( clk , write2_77  , RELUout_F2_2_2  , Final_77_F2_2_2  );
OneRegister RAM_OUT_77_F3_1_1   ( clk , write2_77  , RELUout_F3_1_1  , Final_77_F3_1_1  );
OneRegister RAM_OUT_77_F3_1_2   ( clk , write2_77  , RELUout_F3_1_2  , Final_77_F3_1_2  );
OneRegister RAM_OUT_77_F3_2_1   ( clk , write2_77  , RELUout_F3_2_1  , Final_77_F3_2_1  );
OneRegister RAM_OUT_77_F3_2_2   ( clk , write2_77  , RELUout_F3_2_2  , Final_77_F3_2_2  );
OneRegister RAM_OUT_77_F4_1_1   ( clk , write2_77  , RELUout_F4_1_1  , Final_77_F4_1_1  );
OneRegister RAM_OUT_77_F4_1_2   ( clk , write2_77  , RELUout_F4_1_2  , Final_77_F4_1_2  );
OneRegister RAM_OUT_77_F4_2_1   ( clk , write2_77  , RELUout_F4_2_1  , Final_77_F4_2_1  );
OneRegister RAM_OUT_77_F4_2_2   ( clk , write2_77  , RELUout_F4_2_2  , Final_77_F4_2_2  );
OneRegister RAM_OUT_78_F1_1_1   ( clk , write2_78  , RELUout_F1_1_1  , Final_78_F1_1_1  );
OneRegister RAM_OUT_78_F1_1_2   ( clk , write2_78  , RELUout_F1_1_2  , Final_78_F1_1_2  );
OneRegister RAM_OUT_78_F1_2_1   ( clk , write2_78  , RELUout_F1_2_1  , Final_78_F1_2_1  );
OneRegister RAM_OUT_78_F1_2_2   ( clk , write2_78  , RELUout_F1_2_2  , Final_78_F1_2_2  );
OneRegister RAM_OUT_78_F2_1_1   ( clk , write2_78  , RELUout_F2_1_1  , Final_78_F2_1_1  );
OneRegister RAM_OUT_78_F2_1_2   ( clk , write2_78  , RELUout_F2_1_2  , Final_78_F2_1_2  );
OneRegister RAM_OUT_78_F2_2_1   ( clk , write2_78  , RELUout_F2_2_1  , Final_78_F2_2_1  );
OneRegister RAM_OUT_78_F2_2_2   ( clk , write2_78  , RELUout_F2_2_2  , Final_78_F2_2_2  );
OneRegister RAM_OUT_78_F3_1_1   ( clk , write2_78  , RELUout_F3_1_1  , Final_78_F3_1_1  );
OneRegister RAM_OUT_78_F3_1_2   ( clk , write2_78  , RELUout_F3_1_2  , Final_78_F3_1_2  );
OneRegister RAM_OUT_78_F3_2_1   ( clk , write2_78  , RELUout_F3_2_1  , Final_78_F3_2_1  );
OneRegister RAM_OUT_78_F3_2_2   ( clk , write2_78  , RELUout_F3_2_2  , Final_78_F3_2_2  );
OneRegister RAM_OUT_78_F4_1_1   ( clk , write2_78  , RELUout_F4_1_1  , Final_78_F4_1_1  );
OneRegister RAM_OUT_78_F4_1_2   ( clk , write2_78  , RELUout_F4_1_2  , Final_78_F4_1_2  );
OneRegister RAM_OUT_78_F4_2_1   ( clk , write2_78  , RELUout_F4_2_1  , Final_78_F4_2_1  );
OneRegister RAM_OUT_78_F4_2_2   ( clk , write2_78  , RELUout_F4_2_2  , Final_78_F4_2_2  );
OneRegister RAM_OUT_79_F1_1_1   ( clk , write2_79  , RELUout_F1_1_1  , Final_79_F1_1_1  );
OneRegister RAM_OUT_79_F1_1_2   ( clk , write2_79  , RELUout_F1_1_2  , Final_79_F1_1_2  );
OneRegister RAM_OUT_79_F1_2_1   ( clk , write2_79  , RELUout_F1_2_1  , Final_79_F1_2_1  );
OneRegister RAM_OUT_79_F1_2_2   ( clk , write2_79  , RELUout_F1_2_2  , Final_79_F1_2_2  );
OneRegister RAM_OUT_79_F2_1_1   ( clk , write2_79  , RELUout_F2_1_1  , Final_79_F2_1_1  );
OneRegister RAM_OUT_79_F2_1_2   ( clk , write2_79  , RELUout_F2_1_2  , Final_79_F2_1_2  );
OneRegister RAM_OUT_79_F2_2_1   ( clk , write2_79  , RELUout_F2_2_1  , Final_79_F2_2_1  );
OneRegister RAM_OUT_79_F2_2_2   ( clk , write2_79  , RELUout_F2_2_2  , Final_79_F2_2_2  );
OneRegister RAM_OUT_79_F3_1_1   ( clk , write2_79  , RELUout_F3_1_1  , Final_79_F3_1_1  );
OneRegister RAM_OUT_79_F3_1_2   ( clk , write2_79  , RELUout_F3_1_2  , Final_79_F3_1_2  );
OneRegister RAM_OUT_79_F3_2_1   ( clk , write2_79  , RELUout_F3_2_1  , Final_79_F3_2_1  );
OneRegister RAM_OUT_79_F3_2_2   ( clk , write2_79  , RELUout_F3_2_2  , Final_79_F3_2_2  );
OneRegister RAM_OUT_79_F4_1_1   ( clk , write2_79  , RELUout_F4_1_1  , Final_79_F4_1_1  );
OneRegister RAM_OUT_79_F4_1_2   ( clk , write2_79  , RELUout_F4_1_2  , Final_79_F4_1_2  );
OneRegister RAM_OUT_79_F4_2_1   ( clk , write2_79  , RELUout_F4_2_1  , Final_79_F4_2_1  );
OneRegister RAM_OUT_79_F4_2_2   ( clk , write2_79  , RELUout_F4_2_2  , Final_79_F4_2_2  );
OneRegister RAM_OUT_80_F1_1_1   ( clk , write2_80  , RELUout_F1_1_1  , Final_80_F1_1_1  );
OneRegister RAM_OUT_80_F1_1_2   ( clk , write2_80  , RELUout_F1_1_2  , Final_80_F1_1_2  );
OneRegister RAM_OUT_80_F1_2_1   ( clk , write2_80  , RELUout_F1_2_1  , Final_80_F1_2_1  );
OneRegister RAM_OUT_80_F1_2_2   ( clk , write2_80  , RELUout_F1_2_2  , Final_80_F1_2_2  );
OneRegister RAM_OUT_80_F2_1_1   ( clk , write2_80  , RELUout_F2_1_1  , Final_80_F2_1_1  );
OneRegister RAM_OUT_80_F2_1_2   ( clk , write2_80  , RELUout_F2_1_2  , Final_80_F2_1_2  );
OneRegister RAM_OUT_80_F2_2_1   ( clk , write2_80  , RELUout_F2_2_1  , Final_80_F2_2_1  );
OneRegister RAM_OUT_80_F2_2_2   ( clk , write2_80  , RELUout_F2_2_2  , Final_80_F2_2_2  );
OneRegister RAM_OUT_80_F3_1_1   ( clk , write2_80  , RELUout_F3_1_1  , Final_80_F3_1_1  );
OneRegister RAM_OUT_80_F3_1_2   ( clk , write2_80  , RELUout_F3_1_2  , Final_80_F3_1_2  );
OneRegister RAM_OUT_80_F3_2_1   ( clk , write2_80  , RELUout_F3_2_1  , Final_80_F3_2_1  );
OneRegister RAM_OUT_80_F3_2_2   ( clk , write2_80  , RELUout_F3_2_2  , Final_80_F3_2_2  );
OneRegister RAM_OUT_80_F4_1_1   ( clk , write2_80  , RELUout_F4_1_1  , Final_80_F4_1_1  );
OneRegister RAM_OUT_80_F4_1_2   ( clk , write2_80  , RELUout_F4_1_2  , Final_80_F4_1_2  );
OneRegister RAM_OUT_80_F4_2_1   ( clk , write2_80  , RELUout_F4_2_1  , Final_80_F4_2_1  );
OneRegister RAM_OUT_80_F4_2_2   ( clk , write2_80  , RELUout_F4_2_2  , Final_80_F4_2_2  );
OneRegister RAM_OUT_81_F1_1_1   ( clk , write2_81  , RELUout_F1_1_1  , Final_81_F1_1_1  );
OneRegister RAM_OUT_81_F1_1_2   ( clk , write2_81  , RELUout_F1_1_2  , Final_81_F1_1_2  );
OneRegister RAM_OUT_81_F1_2_1   ( clk , write2_81  , RELUout_F1_2_1  , Final_81_F1_2_1  );
OneRegister RAM_OUT_81_F1_2_2   ( clk , write2_81  , RELUout_F1_2_2  , Final_81_F1_2_2  );
OneRegister RAM_OUT_81_F2_1_1   ( clk , write2_81  , RELUout_F2_1_1  , Final_81_F2_1_1  );
OneRegister RAM_OUT_81_F2_1_2   ( clk , write2_81  , RELUout_F2_1_2  , Final_81_F2_1_2  );
OneRegister RAM_OUT_81_F2_2_1   ( clk , write2_81  , RELUout_F2_2_1  , Final_81_F2_2_1  );
OneRegister RAM_OUT_81_F2_2_2   ( clk , write2_81  , RELUout_F2_2_2  , Final_81_F2_2_2  );
OneRegister RAM_OUT_81_F3_1_1   ( clk , write2_81  , RELUout_F3_1_1  , Final_81_F3_1_1  );
OneRegister RAM_OUT_81_F3_1_2   ( clk , write2_81  , RELUout_F3_1_2  , Final_81_F3_1_2  );
OneRegister RAM_OUT_81_F3_2_1   ( clk , write2_81  , RELUout_F3_2_1  , Final_81_F3_2_1  );
OneRegister RAM_OUT_81_F3_2_2   ( clk , write2_81  , RELUout_F3_2_2  , Final_81_F3_2_2  );
OneRegister RAM_OUT_81_F4_1_1   ( clk , write2_81  , RELUout_F4_1_1  , Final_81_F4_1_1  );
OneRegister RAM_OUT_81_F4_1_2   ( clk , write2_81  , RELUout_F4_1_2  , Final_81_F4_1_2  );
OneRegister RAM_OUT_81_F4_2_1   ( clk , write2_81  , RELUout_F4_2_1  , Final_81_F4_2_1  );
OneRegister RAM_OUT_81_F4_2_2   ( clk , write2_81  , RELUout_F4_2_2  , Final_81_F4_2_2  );
OneRegister RAM_OUT_82_F1_1_1   ( clk , write2_82  , RELUout_F1_1_1  , Final_82_F1_1_1  );
OneRegister RAM_OUT_82_F1_1_2   ( clk , write2_82  , RELUout_F1_1_2  , Final_82_F1_1_2  );
OneRegister RAM_OUT_82_F1_2_1   ( clk , write2_82  , RELUout_F1_2_1  , Final_82_F1_2_1  );
OneRegister RAM_OUT_82_F1_2_2   ( clk , write2_82  , RELUout_F1_2_2  , Final_82_F1_2_2  );
OneRegister RAM_OUT_82_F2_1_1   ( clk , write2_82  , RELUout_F2_1_1  , Final_82_F2_1_1  );
OneRegister RAM_OUT_82_F2_1_2   ( clk , write2_82  , RELUout_F2_1_2  , Final_82_F2_1_2  );
OneRegister RAM_OUT_82_F2_2_1   ( clk , write2_82  , RELUout_F2_2_1  , Final_82_F2_2_1  );
OneRegister RAM_OUT_82_F2_2_2   ( clk , write2_82  , RELUout_F2_2_2  , Final_82_F2_2_2  );
OneRegister RAM_OUT_82_F3_1_1   ( clk , write2_82  , RELUout_F3_1_1  , Final_82_F3_1_1  );
OneRegister RAM_OUT_82_F3_1_2   ( clk , write2_82  , RELUout_F3_1_2  , Final_82_F3_1_2  );
OneRegister RAM_OUT_82_F3_2_1   ( clk , write2_82  , RELUout_F3_2_1  , Final_82_F3_2_1  );
OneRegister RAM_OUT_82_F3_2_2   ( clk , write2_82  , RELUout_F3_2_2  , Final_82_F3_2_2  );
OneRegister RAM_OUT_82_F4_1_1   ( clk , write2_82  , RELUout_F4_1_1  , Final_82_F4_1_1  );
OneRegister RAM_OUT_82_F4_1_2   ( clk , write2_82  , RELUout_F4_1_2  , Final_82_F4_1_2  );
OneRegister RAM_OUT_82_F4_2_1   ( clk , write2_82  , RELUout_F4_2_1  , Final_82_F4_2_1  );
OneRegister RAM_OUT_82_F4_2_2   ( clk , write2_82  , RELUout_F4_2_2  , Final_82_F4_2_2  );
OneRegister RAM_OUT_83_F1_1_1   ( clk , write2_83  , RELUout_F1_1_1  , Final_83_F1_1_1  );
OneRegister RAM_OUT_83_F1_1_2   ( clk , write2_83  , RELUout_F1_1_2  , Final_83_F1_1_2  );
OneRegister RAM_OUT_83_F1_2_1   ( clk , write2_83  , RELUout_F1_2_1  , Final_83_F1_2_1  );
OneRegister RAM_OUT_83_F1_2_2   ( clk , write2_83  , RELUout_F1_2_2  , Final_83_F1_2_2  );
OneRegister RAM_OUT_83_F2_1_1   ( clk , write2_83  , RELUout_F2_1_1  , Final_83_F2_1_1  );
OneRegister RAM_OUT_83_F2_1_2   ( clk , write2_83  , RELUout_F2_1_2  , Final_83_F2_1_2  );
OneRegister RAM_OUT_83_F2_2_1   ( clk , write2_83  , RELUout_F2_2_1  , Final_83_F2_2_1  );
OneRegister RAM_OUT_83_F2_2_2   ( clk , write2_83  , RELUout_F2_2_2  , Final_83_F2_2_2  );
OneRegister RAM_OUT_83_F3_1_1   ( clk , write2_83  , RELUout_F3_1_1  , Final_83_F3_1_1  );
OneRegister RAM_OUT_83_F3_1_2   ( clk , write2_83  , RELUout_F3_1_2  , Final_83_F3_1_2  );
OneRegister RAM_OUT_83_F3_2_1   ( clk , write2_83  , RELUout_F3_2_1  , Final_83_F3_2_1  );
OneRegister RAM_OUT_83_F3_2_2   ( clk , write2_83  , RELUout_F3_2_2  , Final_83_F3_2_2  );
OneRegister RAM_OUT_83_F4_1_1   ( clk , write2_83  , RELUout_F4_1_1  , Final_83_F4_1_1  );
OneRegister RAM_OUT_83_F4_1_2   ( clk , write2_83  , RELUout_F4_1_2  , Final_83_F4_1_2  );
OneRegister RAM_OUT_83_F4_2_1   ( clk , write2_83  , RELUout_F4_2_1  , Final_83_F4_2_1  );
OneRegister RAM_OUT_83_F4_2_2   ( clk , write2_83  , RELUout_F4_2_2  , Final_83_F4_2_2  );
OneRegister RAM_OUT_84_F1_1_1   ( clk , write2_84  , RELUout_F1_1_1  , Final_84_F1_1_1  );
OneRegister RAM_OUT_84_F1_1_2   ( clk , write2_84  , RELUout_F1_1_2  , Final_84_F1_1_2  );
OneRegister RAM_OUT_84_F1_2_1   ( clk , write2_84  , RELUout_F1_2_1  , Final_84_F1_2_1  );
OneRegister RAM_OUT_84_F1_2_2   ( clk , write2_84  , RELUout_F1_2_2  , Final_84_F1_2_2  );
OneRegister RAM_OUT_84_F2_1_1   ( clk , write2_84  , RELUout_F2_1_1  , Final_84_F2_1_1  );
OneRegister RAM_OUT_84_F2_1_2   ( clk , write2_84  , RELUout_F2_1_2  , Final_84_F2_1_2  );
OneRegister RAM_OUT_84_F2_2_1   ( clk , write2_84  , RELUout_F2_2_1  , Final_84_F2_2_1  );
OneRegister RAM_OUT_84_F2_2_2   ( clk , write2_84  , RELUout_F2_2_2  , Final_84_F2_2_2  );
OneRegister RAM_OUT_84_F3_1_1   ( clk , write2_84  , RELUout_F3_1_1  , Final_84_F3_1_1  );
OneRegister RAM_OUT_84_F3_1_2   ( clk , write2_84  , RELUout_F3_1_2  , Final_84_F3_1_2  );
OneRegister RAM_OUT_84_F3_2_1   ( clk , write2_84  , RELUout_F3_2_1  , Final_84_F3_2_1  );
OneRegister RAM_OUT_84_F3_2_2   ( clk , write2_84  , RELUout_F3_2_2  , Final_84_F3_2_2  );
OneRegister RAM_OUT_84_F4_1_1   ( clk , write2_84  , RELUout_F4_1_1  , Final_84_F4_1_1  );
OneRegister RAM_OUT_84_F4_1_2   ( clk , write2_84  , RELUout_F4_1_2  , Final_84_F4_1_2  );
OneRegister RAM_OUT_84_F4_2_1   ( clk , write2_84  , RELUout_F4_2_1  , Final_84_F4_2_1  );
OneRegister RAM_OUT_84_F4_2_2   ( clk , write2_84  , RELUout_F4_2_2  , Final_84_F4_2_2  );
OneRegister RAM_OUT_85_F1_1_1   ( clk , write2_85  , RELUout_F1_1_1  , Final_85_F1_1_1  );
OneRegister RAM_OUT_85_F1_1_2   ( clk , write2_85  , RELUout_F1_1_2  , Final_85_F1_1_2  );
OneRegister RAM_OUT_85_F1_2_1   ( clk , write2_85  , RELUout_F1_2_1  , Final_85_F1_2_1  );
OneRegister RAM_OUT_85_F1_2_2   ( clk , write2_85  , RELUout_F1_2_2  , Final_85_F1_2_2  );
OneRegister RAM_OUT_85_F2_1_1   ( clk , write2_85  , RELUout_F2_1_1  , Final_85_F2_1_1  );
OneRegister RAM_OUT_85_F2_1_2   ( clk , write2_85  , RELUout_F2_1_2  , Final_85_F2_1_2  );
OneRegister RAM_OUT_85_F2_2_1   ( clk , write2_85  , RELUout_F2_2_1  , Final_85_F2_2_1  );
OneRegister RAM_OUT_85_F2_2_2   ( clk , write2_85  , RELUout_F2_2_2  , Final_85_F2_2_2  );
OneRegister RAM_OUT_85_F3_1_1   ( clk , write2_85  , RELUout_F3_1_1  , Final_85_F3_1_1  );
OneRegister RAM_OUT_85_F3_1_2   ( clk , write2_85  , RELUout_F3_1_2  , Final_85_F3_1_2  );
OneRegister RAM_OUT_85_F3_2_1   ( clk , write2_85  , RELUout_F3_2_1  , Final_85_F3_2_1  );
OneRegister RAM_OUT_85_F3_2_2   ( clk , write2_85  , RELUout_F3_2_2  , Final_85_F3_2_2  );
OneRegister RAM_OUT_85_F4_1_1   ( clk , write2_85  , RELUout_F4_1_1  , Final_85_F4_1_1  );
OneRegister RAM_OUT_85_F4_1_2   ( clk , write2_85  , RELUout_F4_1_2  , Final_85_F4_1_2  );
OneRegister RAM_OUT_85_F4_2_1   ( clk , write2_85  , RELUout_F4_2_1  , Final_85_F4_2_1  );
OneRegister RAM_OUT_85_F4_2_2   ( clk , write2_85  , RELUout_F4_2_2  , Final_85_F4_2_2  );
OneRegister RAM_OUT_86_F1_1_1   ( clk , write2_86  , RELUout_F1_1_1  , Final_86_F1_1_1  );
OneRegister RAM_OUT_86_F1_1_2   ( clk , write2_86  , RELUout_F1_1_2  , Final_86_F1_1_2  );
OneRegister RAM_OUT_86_F1_2_1   ( clk , write2_86  , RELUout_F1_2_1  , Final_86_F1_2_1  );
OneRegister RAM_OUT_86_F1_2_2   ( clk , write2_86  , RELUout_F1_2_2  , Final_86_F1_2_2  );
OneRegister RAM_OUT_86_F2_1_1   ( clk , write2_86  , RELUout_F2_1_1  , Final_86_F2_1_1  );
OneRegister RAM_OUT_86_F2_1_2   ( clk , write2_86  , RELUout_F2_1_2  , Final_86_F2_1_2  );
OneRegister RAM_OUT_86_F2_2_1   ( clk , write2_86  , RELUout_F2_2_1  , Final_86_F2_2_1  );
OneRegister RAM_OUT_86_F2_2_2   ( clk , write2_86  , RELUout_F2_2_2  , Final_86_F2_2_2  );
OneRegister RAM_OUT_86_F3_1_1   ( clk , write2_86  , RELUout_F3_1_1  , Final_86_F3_1_1  );
OneRegister RAM_OUT_86_F3_1_2   ( clk , write2_86  , RELUout_F3_1_2  , Final_86_F3_1_2  );
OneRegister RAM_OUT_86_F3_2_1   ( clk , write2_86  , RELUout_F3_2_1  , Final_86_F3_2_1  );
OneRegister RAM_OUT_86_F3_2_2   ( clk , write2_86  , RELUout_F3_2_2  , Final_86_F3_2_2  );
OneRegister RAM_OUT_86_F4_1_1   ( clk , write2_86  , RELUout_F4_1_1  , Final_86_F4_1_1  );
OneRegister RAM_OUT_86_F4_1_2   ( clk , write2_86  , RELUout_F4_1_2  , Final_86_F4_1_2  );
OneRegister RAM_OUT_86_F4_2_1   ( clk , write2_86  , RELUout_F4_2_1  , Final_86_F4_2_1  );
OneRegister RAM_OUT_86_F4_2_2   ( clk , write2_86  , RELUout_F4_2_2  , Final_86_F4_2_2  );
OneRegister RAM_OUT_87_F1_1_1   ( clk , write2_87  , RELUout_F1_1_1  , Final_87_F1_1_1  );
OneRegister RAM_OUT_87_F1_1_2   ( clk , write2_87  , RELUout_F1_1_2  , Final_87_F1_1_2  );
OneRegister RAM_OUT_87_F1_2_1   ( clk , write2_87  , RELUout_F1_2_1  , Final_87_F1_2_1  );
OneRegister RAM_OUT_87_F1_2_2   ( clk , write2_87  , RELUout_F1_2_2  , Final_87_F1_2_2  );
OneRegister RAM_OUT_87_F2_1_1   ( clk , write2_87  , RELUout_F2_1_1  , Final_87_F2_1_1  );
OneRegister RAM_OUT_87_F2_1_2   ( clk , write2_87  , RELUout_F2_1_2  , Final_87_F2_1_2  );
OneRegister RAM_OUT_87_F2_2_1   ( clk , write2_87  , RELUout_F2_2_1  , Final_87_F2_2_1  );
OneRegister RAM_OUT_87_F2_2_2   ( clk , write2_87  , RELUout_F2_2_2  , Final_87_F2_2_2  );
OneRegister RAM_OUT_87_F3_1_1   ( clk , write2_87  , RELUout_F3_1_1  , Final_87_F3_1_1  );
OneRegister RAM_OUT_87_F3_1_2   ( clk , write2_87  , RELUout_F3_1_2  , Final_87_F3_1_2  );
OneRegister RAM_OUT_87_F3_2_1   ( clk , write2_87  , RELUout_F3_2_1  , Final_87_F3_2_1  );
OneRegister RAM_OUT_87_F3_2_2   ( clk , write2_87  , RELUout_F3_2_2  , Final_87_F3_2_2  );
OneRegister RAM_OUT_87_F4_1_1   ( clk , write2_87  , RELUout_F4_1_1  , Final_87_F4_1_1  );
OneRegister RAM_OUT_87_F4_1_2   ( clk , write2_87  , RELUout_F4_1_2  , Final_87_F4_1_2  );
OneRegister RAM_OUT_87_F4_2_1   ( clk , write2_87  , RELUout_F4_2_1  , Final_87_F4_2_1  );
OneRegister RAM_OUT_87_F4_2_2   ( clk , write2_87  , RELUout_F4_2_2  , Final_87_F4_2_2  );
OneRegister RAM_OUT_88_F1_1_1   ( clk , write2_88  , RELUout_F1_1_1  , Final_88_F1_1_1  );
OneRegister RAM_OUT_88_F1_1_2   ( clk , write2_88  , RELUout_F1_1_2  , Final_88_F1_1_2  );
OneRegister RAM_OUT_88_F1_2_1   ( clk , write2_88  , RELUout_F1_2_1  , Final_88_F1_2_1  );
OneRegister RAM_OUT_88_F1_2_2   ( clk , write2_88  , RELUout_F1_2_2  , Final_88_F1_2_2  );
OneRegister RAM_OUT_88_F2_1_1   ( clk , write2_88  , RELUout_F2_1_1  , Final_88_F2_1_1  );
OneRegister RAM_OUT_88_F2_1_2   ( clk , write2_88  , RELUout_F2_1_2  , Final_88_F2_1_2  );
OneRegister RAM_OUT_88_F2_2_1   ( clk , write2_88  , RELUout_F2_2_1  , Final_88_F2_2_1  );
OneRegister RAM_OUT_88_F2_2_2   ( clk , write2_88  , RELUout_F2_2_2  , Final_88_F2_2_2  );
OneRegister RAM_OUT_88_F3_1_1   ( clk , write2_88  , RELUout_F3_1_1  , Final_88_F3_1_1  );
OneRegister RAM_OUT_88_F3_1_2   ( clk , write2_88  , RELUout_F3_1_2  , Final_88_F3_1_2  );
OneRegister RAM_OUT_88_F3_2_1   ( clk , write2_88  , RELUout_F3_2_1  , Final_88_F3_2_1  );
OneRegister RAM_OUT_88_F3_2_2   ( clk , write2_88  , RELUout_F3_2_2  , Final_88_F3_2_2  );
OneRegister RAM_OUT_88_F4_1_1   ( clk , write2_88  , RELUout_F4_1_1  , Final_88_F4_1_1  );
OneRegister RAM_OUT_88_F4_1_2   ( clk , write2_88  , RELUout_F4_1_2  , Final_88_F4_1_2  );
OneRegister RAM_OUT_88_F4_2_1   ( clk , write2_88  , RELUout_F4_2_1  , Final_88_F4_2_1  );
OneRegister RAM_OUT_88_F4_2_2   ( clk , write2_88  , RELUout_F4_2_2  , Final_88_F4_2_2  );
OneRegister RAM_OUT_89_F1_1_1   ( clk , write2_89  , RELUout_F1_1_1  , Final_89_F1_1_1  );
OneRegister RAM_OUT_89_F1_1_2   ( clk , write2_89  , RELUout_F1_1_2  , Final_89_F1_1_2  );
OneRegister RAM_OUT_89_F1_2_1   ( clk , write2_89  , RELUout_F1_2_1  , Final_89_F1_2_1  );
OneRegister RAM_OUT_89_F1_2_2   ( clk , write2_89  , RELUout_F1_2_2  , Final_89_F1_2_2  );
OneRegister RAM_OUT_89_F2_1_1   ( clk , write2_89  , RELUout_F2_1_1  , Final_89_F2_1_1  );
OneRegister RAM_OUT_89_F2_1_2   ( clk , write2_89  , RELUout_F2_1_2  , Final_89_F2_1_2  );
OneRegister RAM_OUT_89_F2_2_1   ( clk , write2_89  , RELUout_F2_2_1  , Final_89_F2_2_1  );
OneRegister RAM_OUT_89_F2_2_2   ( clk , write2_89  , RELUout_F2_2_2  , Final_89_F2_2_2  );
OneRegister RAM_OUT_89_F3_1_1   ( clk , write2_89  , RELUout_F3_1_1  , Final_89_F3_1_1  );
OneRegister RAM_OUT_89_F3_1_2   ( clk , write2_89  , RELUout_F3_1_2  , Final_89_F3_1_2  );
OneRegister RAM_OUT_89_F3_2_1   ( clk , write2_89  , RELUout_F3_2_1  , Final_89_F3_2_1  );
OneRegister RAM_OUT_89_F3_2_2   ( clk , write2_89  , RELUout_F3_2_2  , Final_89_F3_2_2  );
OneRegister RAM_OUT_89_F4_1_1   ( clk , write2_89  , RELUout_F4_1_1  , Final_89_F4_1_1  );
OneRegister RAM_OUT_89_F4_1_2   ( clk , write2_89  , RELUout_F4_1_2  , Final_89_F4_1_2  );
OneRegister RAM_OUT_89_F4_2_1   ( clk , write2_89  , RELUout_F4_2_1  , Final_89_F4_2_1  );
OneRegister RAM_OUT_89_F4_2_2   ( clk , write2_89  , RELUout_F4_2_2  , Final_89_F4_2_2  );
OneRegister RAM_OUT_90_F1_1_1   ( clk , write2_90  , RELUout_F1_1_1  , Final_90_F1_1_1  );
OneRegister RAM_OUT_90_F1_1_2   ( clk , write2_90  , RELUout_F1_1_2  , Final_90_F1_1_2  );
OneRegister RAM_OUT_90_F1_2_1   ( clk , write2_90  , RELUout_F1_2_1  , Final_90_F1_2_1  );
OneRegister RAM_OUT_90_F1_2_2   ( clk , write2_90  , RELUout_F1_2_2  , Final_90_F1_2_2  );
OneRegister RAM_OUT_90_F2_1_1   ( clk , write2_90  , RELUout_F2_1_1  , Final_90_F2_1_1  );
OneRegister RAM_OUT_90_F2_1_2   ( clk , write2_90  , RELUout_F2_1_2  , Final_90_F2_1_2  );
OneRegister RAM_OUT_90_F2_2_1   ( clk , write2_90  , RELUout_F2_2_1  , Final_90_F2_2_1  );
OneRegister RAM_OUT_90_F2_2_2   ( clk , write2_90  , RELUout_F2_2_2  , Final_90_F2_2_2  );
OneRegister RAM_OUT_90_F3_1_1   ( clk , write2_90  , RELUout_F3_1_1  , Final_90_F3_1_1  );
OneRegister RAM_OUT_90_F3_1_2   ( clk , write2_90  , RELUout_F3_1_2  , Final_90_F3_1_2  );
OneRegister RAM_OUT_90_F3_2_1   ( clk , write2_90  , RELUout_F3_2_1  , Final_90_F3_2_1  );
OneRegister RAM_OUT_90_F3_2_2   ( clk , write2_90  , RELUout_F3_2_2  , Final_90_F3_2_2  );
OneRegister RAM_OUT_90_F4_1_1   ( clk , write2_90  , RELUout_F4_1_1  , Final_90_F4_1_1  );
OneRegister RAM_OUT_90_F4_1_2   ( clk , write2_90  , RELUout_F4_1_2  , Final_90_F4_1_2  );
OneRegister RAM_OUT_90_F4_2_1   ( clk , write2_90  , RELUout_F4_2_1  , Final_90_F4_2_1  );
OneRegister RAM_OUT_90_F4_2_2   ( clk , write2_90  , RELUout_F4_2_2  , Final_90_F4_2_2  );
OneRegister RAM_OUT_91_F1_1_1   ( clk , write2_91  , RELUout_F1_1_1  , Final_91_F1_1_1  );
OneRegister RAM_OUT_91_F1_1_2   ( clk , write2_91  , RELUout_F1_1_2  , Final_91_F1_1_2  );
OneRegister RAM_OUT_91_F1_2_1   ( clk , write2_91  , RELUout_F1_2_1  , Final_91_F1_2_1  );
OneRegister RAM_OUT_91_F1_2_2   ( clk , write2_91  , RELUout_F1_2_2  , Final_91_F1_2_2  );
OneRegister RAM_OUT_91_F2_1_1   ( clk , write2_91  , RELUout_F2_1_1  , Final_91_F2_1_1  );
OneRegister RAM_OUT_91_F2_1_2   ( clk , write2_91  , RELUout_F2_1_2  , Final_91_F2_1_2  );
OneRegister RAM_OUT_91_F2_2_1   ( clk , write2_91  , RELUout_F2_2_1  , Final_91_F2_2_1  );
OneRegister RAM_OUT_91_F2_2_2   ( clk , write2_91  , RELUout_F2_2_2  , Final_91_F2_2_2  );
OneRegister RAM_OUT_91_F3_1_1   ( clk , write2_91  , RELUout_F3_1_1  , Final_91_F3_1_1  );
OneRegister RAM_OUT_91_F3_1_2   ( clk , write2_91  , RELUout_F3_1_2  , Final_91_F3_1_2  );
OneRegister RAM_OUT_91_F3_2_1   ( clk , write2_91  , RELUout_F3_2_1  , Final_91_F3_2_1  );
OneRegister RAM_OUT_91_F3_2_2   ( clk , write2_91  , RELUout_F3_2_2  , Final_91_F3_2_2  );
OneRegister RAM_OUT_91_F4_1_1   ( clk , write2_91  , RELUout_F4_1_1  , Final_91_F4_1_1  );
OneRegister RAM_OUT_91_F4_1_2   ( clk , write2_91  , RELUout_F4_1_2  , Final_91_F4_1_2  );
OneRegister RAM_OUT_91_F4_2_1   ( clk , write2_91  , RELUout_F4_2_1  , Final_91_F4_2_1  );
OneRegister RAM_OUT_91_F4_2_2   ( clk , write2_91  , RELUout_F4_2_2  , Final_91_F4_2_2  );
OneRegister RAM_OUT_92_F1_1_1   ( clk , write2_92  , RELUout_F1_1_1  , Final_92_F1_1_1  );
OneRegister RAM_OUT_92_F1_1_2   ( clk , write2_92  , RELUout_F1_1_2  , Final_92_F1_1_2  );
OneRegister RAM_OUT_92_F1_2_1   ( clk , write2_92  , RELUout_F1_2_1  , Final_92_F1_2_1  );
OneRegister RAM_OUT_92_F1_2_2   ( clk , write2_92  , RELUout_F1_2_2  , Final_92_F1_2_2  );
OneRegister RAM_OUT_92_F2_1_1   ( clk , write2_92  , RELUout_F2_1_1  , Final_92_F2_1_1  );
OneRegister RAM_OUT_92_F2_1_2   ( clk , write2_92  , RELUout_F2_1_2  , Final_92_F2_1_2  );
OneRegister RAM_OUT_92_F2_2_1   ( clk , write2_92  , RELUout_F2_2_1  , Final_92_F2_2_1  );
OneRegister RAM_OUT_92_F2_2_2   ( clk , write2_92  , RELUout_F2_2_2  , Final_92_F2_2_2  );
OneRegister RAM_OUT_92_F3_1_1   ( clk , write2_92  , RELUout_F3_1_1  , Final_92_F3_1_1  );
OneRegister RAM_OUT_92_F3_1_2   ( clk , write2_92  , RELUout_F3_1_2  , Final_92_F3_1_2  );
OneRegister RAM_OUT_92_F3_2_1   ( clk , write2_92  , RELUout_F3_2_1  , Final_92_F3_2_1  );
OneRegister RAM_OUT_92_F3_2_2   ( clk , write2_92  , RELUout_F3_2_2  , Final_92_F3_2_2  );
OneRegister RAM_OUT_92_F4_1_1   ( clk , write2_92  , RELUout_F4_1_1  , Final_92_F4_1_1  );
OneRegister RAM_OUT_92_F4_1_2   ( clk , write2_92  , RELUout_F4_1_2  , Final_92_F4_1_2  );
OneRegister RAM_OUT_92_F4_2_1   ( clk , write2_92  , RELUout_F4_2_1  , Final_92_F4_2_1  );
OneRegister RAM_OUT_92_F4_2_2   ( clk , write2_92  , RELUout_F4_2_2  , Final_92_F4_2_2  );
OneRegister RAM_OUT_93_F1_1_1   ( clk , write2_93  , RELUout_F1_1_1  , Final_93_F1_1_1  );
OneRegister RAM_OUT_93_F1_1_2   ( clk , write2_93  , RELUout_F1_1_2  , Final_93_F1_1_2  );
OneRegister RAM_OUT_93_F1_2_1   ( clk , write2_93  , RELUout_F1_2_1  , Final_93_F1_2_1  );
OneRegister RAM_OUT_93_F1_2_2   ( clk , write2_93  , RELUout_F1_2_2  , Final_93_F1_2_2  );
OneRegister RAM_OUT_93_F2_1_1   ( clk , write2_93  , RELUout_F2_1_1  , Final_93_F2_1_1  );
OneRegister RAM_OUT_93_F2_1_2   ( clk , write2_93  , RELUout_F2_1_2  , Final_93_F2_1_2  );
OneRegister RAM_OUT_93_F2_2_1   ( clk , write2_93  , RELUout_F2_2_1  , Final_93_F2_2_1  );
OneRegister RAM_OUT_93_F2_2_2   ( clk , write2_93  , RELUout_F2_2_2  , Final_93_F2_2_2  );
OneRegister RAM_OUT_93_F3_1_1   ( clk , write2_93  , RELUout_F3_1_1  , Final_93_F3_1_1  );
OneRegister RAM_OUT_93_F3_1_2   ( clk , write2_93  , RELUout_F3_1_2  , Final_93_F3_1_2  );
OneRegister RAM_OUT_93_F3_2_1   ( clk , write2_93  , RELUout_F3_2_1  , Final_93_F3_2_1  );
OneRegister RAM_OUT_93_F3_2_2   ( clk , write2_93  , RELUout_F3_2_2  , Final_93_F3_2_2  );
OneRegister RAM_OUT_93_F4_1_1   ( clk , write2_93  , RELUout_F4_1_1  , Final_93_F4_1_1  );
OneRegister RAM_OUT_93_F4_1_2   ( clk , write2_93  , RELUout_F4_1_2  , Final_93_F4_1_2  );
OneRegister RAM_OUT_93_F4_2_1   ( clk , write2_93  , RELUout_F4_2_1  , Final_93_F4_2_1  );
OneRegister RAM_OUT_93_F4_2_2   ( clk , write2_93  , RELUout_F4_2_2  , Final_93_F4_2_2  );
OneRegister RAM_OUT_94_F1_1_1   ( clk , write2_94  , RELUout_F1_1_1  , Final_94_F1_1_1  );
OneRegister RAM_OUT_94_F1_1_2   ( clk , write2_94  , RELUout_F1_1_2  , Final_94_F1_1_2  );
OneRegister RAM_OUT_94_F1_2_1   ( clk , write2_94  , RELUout_F1_2_1  , Final_94_F1_2_1  );
OneRegister RAM_OUT_94_F1_2_2   ( clk , write2_94  , RELUout_F1_2_2  , Final_94_F1_2_2  );
OneRegister RAM_OUT_94_F2_1_1   ( clk , write2_94  , RELUout_F2_1_1  , Final_94_F2_1_1  );
OneRegister RAM_OUT_94_F2_1_2   ( clk , write2_94  , RELUout_F2_1_2  , Final_94_F2_1_2  );
OneRegister RAM_OUT_94_F2_2_1   ( clk , write2_94  , RELUout_F2_2_1  , Final_94_F2_2_1  );
OneRegister RAM_OUT_94_F2_2_2   ( clk , write2_94  , RELUout_F2_2_2  , Final_94_F2_2_2  );
OneRegister RAM_OUT_94_F3_1_1   ( clk , write2_94  , RELUout_F3_1_1  , Final_94_F3_1_1  );
OneRegister RAM_OUT_94_F3_1_2   ( clk , write2_94  , RELUout_F3_1_2  , Final_94_F3_1_2  );
OneRegister RAM_OUT_94_F3_2_1   ( clk , write2_94  , RELUout_F3_2_1  , Final_94_F3_2_1  );
OneRegister RAM_OUT_94_F3_2_2   ( clk , write2_94  , RELUout_F3_2_2  , Final_94_F3_2_2  );
OneRegister RAM_OUT_94_F4_1_1   ( clk , write2_94  , RELUout_F4_1_1  , Final_94_F4_1_1  );
OneRegister RAM_OUT_94_F4_1_2   ( clk , write2_94  , RELUout_F4_1_2  , Final_94_F4_1_2  );
OneRegister RAM_OUT_94_F4_2_1   ( clk , write2_94  , RELUout_F4_2_1  , Final_94_F4_2_1  );
OneRegister RAM_OUT_94_F4_2_2   ( clk , write2_94  , RELUout_F4_2_2  , Final_94_F4_2_2  );
OneRegister RAM_OUT_95_F1_1_1   ( clk , write2_95  , RELUout_F1_1_1  , Final_95_F1_1_1  );
OneRegister RAM_OUT_95_F1_1_2   ( clk , write2_95  , RELUout_F1_1_2  , Final_95_F1_1_2  );
OneRegister RAM_OUT_95_F1_2_1   ( clk , write2_95  , RELUout_F1_2_1  , Final_95_F1_2_1  );
OneRegister RAM_OUT_95_F1_2_2   ( clk , write2_95  , RELUout_F1_2_2  , Final_95_F1_2_2  );
OneRegister RAM_OUT_95_F2_1_1   ( clk , write2_95  , RELUout_F2_1_1  , Final_95_F2_1_1  );
OneRegister RAM_OUT_95_F2_1_2   ( clk , write2_95  , RELUout_F2_1_2  , Final_95_F2_1_2  );
OneRegister RAM_OUT_95_F2_2_1   ( clk , write2_95  , RELUout_F2_2_1  , Final_95_F2_2_1  );
OneRegister RAM_OUT_95_F2_2_2   ( clk , write2_95  , RELUout_F2_2_2  , Final_95_F2_2_2  );
OneRegister RAM_OUT_95_F3_1_1   ( clk , write2_95  , RELUout_F3_1_1  , Final_95_F3_1_1  );
OneRegister RAM_OUT_95_F3_1_2   ( clk , write2_95  , RELUout_F3_1_2  , Final_95_F3_1_2  );
OneRegister RAM_OUT_95_F3_2_1   ( clk , write2_95  , RELUout_F3_2_1  , Final_95_F3_2_1  );
OneRegister RAM_OUT_95_F3_2_2   ( clk , write2_95  , RELUout_F3_2_2  , Final_95_F3_2_2  );
OneRegister RAM_OUT_95_F4_1_1   ( clk , write2_95  , RELUout_F4_1_1  , Final_95_F4_1_1  );
OneRegister RAM_OUT_95_F4_1_2   ( clk , write2_95  , RELUout_F4_1_2  , Final_95_F4_1_2  );
OneRegister RAM_OUT_95_F4_2_1   ( clk , write2_95  , RELUout_F4_2_1  , Final_95_F4_2_1  );
OneRegister RAM_OUT_95_F4_2_2   ( clk , write2_95  , RELUout_F4_2_2  , Final_95_F4_2_2  );
OneRegister RAM_OUT_96_F1_1_1   ( clk , write2_96  , RELUout_F1_1_1  , Final_96_F1_1_1  );
OneRegister RAM_OUT_96_F1_1_2   ( clk , write2_96  , RELUout_F1_1_2  , Final_96_F1_1_2  );
OneRegister RAM_OUT_96_F1_2_1   ( clk , write2_96  , RELUout_F1_2_1  , Final_96_F1_2_1  );
OneRegister RAM_OUT_96_F1_2_2   ( clk , write2_96  , RELUout_F1_2_2  , Final_96_F1_2_2  );
OneRegister RAM_OUT_96_F2_1_1   ( clk , write2_96  , RELUout_F2_1_1  , Final_96_F2_1_1  );
OneRegister RAM_OUT_96_F2_1_2   ( clk , write2_96  , RELUout_F2_1_2  , Final_96_F2_1_2  );
OneRegister RAM_OUT_96_F2_2_1   ( clk , write2_96  , RELUout_F2_2_1  , Final_96_F2_2_1  );
OneRegister RAM_OUT_96_F2_2_2   ( clk , write2_96  , RELUout_F2_2_2  , Final_96_F2_2_2  );
OneRegister RAM_OUT_96_F3_1_1   ( clk , write2_96  , RELUout_F3_1_1  , Final_96_F3_1_1  );
OneRegister RAM_OUT_96_F3_1_2   ( clk , write2_96  , RELUout_F3_1_2  , Final_96_F3_1_2  );
OneRegister RAM_OUT_96_F3_2_1   ( clk , write2_96  , RELUout_F3_2_1  , Final_96_F3_2_1  );
OneRegister RAM_OUT_96_F3_2_2   ( clk , write2_96  , RELUout_F3_2_2  , Final_96_F3_2_2  );
OneRegister RAM_OUT_96_F4_1_1   ( clk , write2_96  , RELUout_F4_1_1  , Final_96_F4_1_1  );
OneRegister RAM_OUT_96_F4_1_2   ( clk , write2_96  , RELUout_F4_1_2  , Final_96_F4_1_2  );
OneRegister RAM_OUT_96_F4_2_1   ( clk , write2_96  , RELUout_F4_2_1  , Final_96_F4_2_1  );
OneRegister RAM_OUT_96_F4_2_2   ( clk , write2_96  , RELUout_F4_2_2  , Final_96_F4_2_2  );
OneRegister RAM_OUT_97_F1_1_1   ( clk , write2_97  , RELUout_F1_1_1  , Final_97_F1_1_1  );
OneRegister RAM_OUT_97_F1_1_2   ( clk , write2_97  , RELUout_F1_1_2  , Final_97_F1_1_2  );
OneRegister RAM_OUT_97_F1_2_1   ( clk , write2_97  , RELUout_F1_2_1  , Final_97_F1_2_1  );
OneRegister RAM_OUT_97_F1_2_2   ( clk , write2_97  , RELUout_F1_2_2  , Final_97_F1_2_2  );
OneRegister RAM_OUT_97_F2_1_1   ( clk , write2_97  , RELUout_F2_1_1  , Final_97_F2_1_1  );
OneRegister RAM_OUT_97_F2_1_2   ( clk , write2_97  , RELUout_F2_1_2  , Final_97_F2_1_2  );
OneRegister RAM_OUT_97_F2_2_1   ( clk , write2_97  , RELUout_F2_2_1  , Final_97_F2_2_1  );
OneRegister RAM_OUT_97_F2_2_2   ( clk , write2_97  , RELUout_F2_2_2  , Final_97_F2_2_2  );
OneRegister RAM_OUT_97_F3_1_1   ( clk , write2_97  , RELUout_F3_1_1  , Final_97_F3_1_1  );
OneRegister RAM_OUT_97_F3_1_2   ( clk , write2_97  , RELUout_F3_1_2  , Final_97_F3_1_2  );
OneRegister RAM_OUT_97_F3_2_1   ( clk , write2_97  , RELUout_F3_2_1  , Final_97_F3_2_1  );
OneRegister RAM_OUT_97_F3_2_2   ( clk , write2_97  , RELUout_F3_2_2  , Final_97_F3_2_2  );
OneRegister RAM_OUT_97_F4_1_1   ( clk , write2_97  , RELUout_F4_1_1  , Final_97_F4_1_1  );
OneRegister RAM_OUT_97_F4_1_2   ( clk , write2_97  , RELUout_F4_1_2  , Final_97_F4_1_2  );
OneRegister RAM_OUT_97_F4_2_1   ( clk , write2_97  , RELUout_F4_2_1  , Final_97_F4_2_1  );
OneRegister RAM_OUT_97_F4_2_2   ( clk , write2_97  , RELUout_F4_2_2  , Final_97_F4_2_2  );
OneRegister RAM_OUT_98_F1_1_1   ( clk , write2_98  , RELUout_F1_1_1  , Final_98_F1_1_1  );
OneRegister RAM_OUT_98_F1_1_2   ( clk , write2_98  , RELUout_F1_1_2  , Final_98_F1_1_2  );
OneRegister RAM_OUT_98_F1_2_1   ( clk , write2_98  , RELUout_F1_2_1  , Final_98_F1_2_1  );
OneRegister RAM_OUT_98_F1_2_2   ( clk , write2_98  , RELUout_F1_2_2  , Final_98_F1_2_2  );
OneRegister RAM_OUT_98_F2_1_1   ( clk , write2_98  , RELUout_F2_1_1  , Final_98_F2_1_1  );
OneRegister RAM_OUT_98_F2_1_2   ( clk , write2_98  , RELUout_F2_1_2  , Final_98_F2_1_2  );
OneRegister RAM_OUT_98_F2_2_1   ( clk , write2_98  , RELUout_F2_2_1  , Final_98_F2_2_1  );
OneRegister RAM_OUT_98_F2_2_2   ( clk , write2_98  , RELUout_F2_2_2  , Final_98_F2_2_2  );
OneRegister RAM_OUT_98_F3_1_1   ( clk , write2_98  , RELUout_F3_1_1  , Final_98_F3_1_1  );
OneRegister RAM_OUT_98_F3_1_2   ( clk , write2_98  , RELUout_F3_1_2  , Final_98_F3_1_2  );
OneRegister RAM_OUT_98_F3_2_1   ( clk , write2_98  , RELUout_F3_2_1  , Final_98_F3_2_1  );
OneRegister RAM_OUT_98_F3_2_2   ( clk , write2_98  , RELUout_F3_2_2  , Final_98_F3_2_2  );
OneRegister RAM_OUT_98_F4_1_1   ( clk , write2_98  , RELUout_F4_1_1  , Final_98_F4_1_1  );
OneRegister RAM_OUT_98_F4_1_2   ( clk , write2_98  , RELUout_F4_1_2  , Final_98_F4_1_2  );
OneRegister RAM_OUT_98_F4_2_1   ( clk , write2_98  , RELUout_F4_2_1  , Final_98_F4_2_1  );
OneRegister RAM_OUT_98_F4_2_2   ( clk , write2_98  , RELUout_F4_2_2  , Final_98_F4_2_2  );
OneRegister RAM_OUT_99_F1_1_1   ( clk , write2_99  , RELUout_F1_1_1  , Final_99_F1_1_1  );
OneRegister RAM_OUT_99_F1_1_2   ( clk , write2_99  , RELUout_F1_1_2  , Final_99_F1_1_2  );
OneRegister RAM_OUT_99_F1_2_1   ( clk , write2_99  , RELUout_F1_2_1  , Final_99_F1_2_1  );
OneRegister RAM_OUT_99_F1_2_2   ( clk , write2_99  , RELUout_F1_2_2  , Final_99_F1_2_2  );
OneRegister RAM_OUT_99_F2_1_1   ( clk , write2_99  , RELUout_F2_1_1  , Final_99_F2_1_1  );
OneRegister RAM_OUT_99_F2_1_2   ( clk , write2_99  , RELUout_F2_1_2  , Final_99_F2_1_2  );
OneRegister RAM_OUT_99_F2_2_1   ( clk , write2_99  , RELUout_F2_2_1  , Final_99_F2_2_1  );
OneRegister RAM_OUT_99_F2_2_2   ( clk , write2_99  , RELUout_F2_2_2  , Final_99_F2_2_2  );
OneRegister RAM_OUT_99_F3_1_1   ( clk , write2_99  , RELUout_F3_1_1  , Final_99_F3_1_1  );
OneRegister RAM_OUT_99_F3_1_2   ( clk , write2_99  , RELUout_F3_1_2  , Final_99_F3_1_2  );
OneRegister RAM_OUT_99_F3_2_1   ( clk , write2_99  , RELUout_F3_2_1  , Final_99_F3_2_1  );
OneRegister RAM_OUT_99_F3_2_2   ( clk , write2_99  , RELUout_F3_2_2  , Final_99_F3_2_2  );
OneRegister RAM_OUT_99_F4_1_1   ( clk , write2_99  , RELUout_F4_1_1  , Final_99_F4_1_1  );
OneRegister RAM_OUT_99_F4_1_2   ( clk , write2_99  , RELUout_F4_1_2  , Final_99_F4_1_2  );
OneRegister RAM_OUT_99_F4_2_1   ( clk , write2_99  , RELUout_F4_2_1  , Final_99_F4_2_1  );
OneRegister RAM_OUT_99_F4_2_2   ( clk , write2_99  , RELUout_F4_2_2  , Final_99_F4_2_2  );
OneRegister RAM_OUT_100_F1_1_1   ( clk , write2_100  , RELUout_F1_1_1  , Final_100_F1_1_1  );
OneRegister RAM_OUT_100_F1_1_2   ( clk , write2_100  , RELUout_F1_1_2  , Final_100_F1_1_2  );
OneRegister RAM_OUT_100_F1_2_1   ( clk , write2_100  , RELUout_F1_2_1  , Final_100_F1_2_1  );
OneRegister RAM_OUT_100_F1_2_2   ( clk , write2_100  , RELUout_F1_2_2  , Final_100_F1_2_2  );
OneRegister RAM_OUT_100_F2_1_1   ( clk , write2_100  , RELUout_F2_1_1  , Final_100_F2_1_1  );
OneRegister RAM_OUT_100_F2_1_2   ( clk , write2_100  , RELUout_F2_1_2  , Final_100_F2_1_2  );
OneRegister RAM_OUT_100_F2_2_1   ( clk , write2_100  , RELUout_F2_2_1  , Final_100_F2_2_1  );
OneRegister RAM_OUT_100_F2_2_2   ( clk , write2_100  , RELUout_F2_2_2  , Final_100_F2_2_2  );
OneRegister RAM_OUT_100_F3_1_1   ( clk , write2_100  , RELUout_F3_1_1  , Final_100_F3_1_1  );
OneRegister RAM_OUT_100_F3_1_2   ( clk , write2_100  , RELUout_F3_1_2  , Final_100_F3_1_2  );
OneRegister RAM_OUT_100_F3_2_1   ( clk , write2_100  , RELUout_F3_2_1  , Final_100_F3_2_1  );
OneRegister RAM_OUT_100_F3_2_2   ( clk , write2_100  , RELUout_F3_2_2  , Final_100_F3_2_2  );
OneRegister RAM_OUT_100_F4_1_1   ( clk , write2_100  , RELUout_F4_1_1  , Final_100_F4_1_1  );
OneRegister RAM_OUT_100_F4_1_2   ( clk , write2_100  , RELUout_F4_1_2  , Final_100_F4_1_2  );
OneRegister RAM_OUT_100_F4_2_1   ( clk , write2_100  , RELUout_F4_2_1  , Final_100_F4_2_1  );
OneRegister RAM_OUT_100_F4_2_2   ( clk , write2_100  , RELUout_F4_2_2  , Final_100_F4_2_2  );
OneRegister RAM_OUT_101_F1_1_1   ( clk , write2_101  , RELUout_F1_1_1  , Final_101_F1_1_1  );
OneRegister RAM_OUT_101_F1_1_2   ( clk , write2_101  , RELUout_F1_1_2  , Final_101_F1_1_2  );
OneRegister RAM_OUT_101_F1_2_1   ( clk , write2_101  , RELUout_F1_2_1  , Final_101_F1_2_1  );
OneRegister RAM_OUT_101_F1_2_2   ( clk , write2_101  , RELUout_F1_2_2  , Final_101_F1_2_2  );
OneRegister RAM_OUT_101_F2_1_1   ( clk , write2_101  , RELUout_F2_1_1  , Final_101_F2_1_1  );
OneRegister RAM_OUT_101_F2_1_2   ( clk , write2_101  , RELUout_F2_1_2  , Final_101_F2_1_2  );
OneRegister RAM_OUT_101_F2_2_1   ( clk , write2_101  , RELUout_F2_2_1  , Final_101_F2_2_1  );
OneRegister RAM_OUT_101_F2_2_2   ( clk , write2_101  , RELUout_F2_2_2  , Final_101_F2_2_2  );
OneRegister RAM_OUT_101_F3_1_1   ( clk , write2_101  , RELUout_F3_1_1  , Final_101_F3_1_1  );
OneRegister RAM_OUT_101_F3_1_2   ( clk , write2_101  , RELUout_F3_1_2  , Final_101_F3_1_2  );
OneRegister RAM_OUT_101_F3_2_1   ( clk , write2_101  , RELUout_F3_2_1  , Final_101_F3_2_1  );
OneRegister RAM_OUT_101_F3_2_2   ( clk , write2_101  , RELUout_F3_2_2  , Final_101_F3_2_2  );
OneRegister RAM_OUT_101_F4_1_1   ( clk , write2_101  , RELUout_F4_1_1  , Final_101_F4_1_1  );
OneRegister RAM_OUT_101_F4_1_2   ( clk , write2_101  , RELUout_F4_1_2  , Final_101_F4_1_2  );
OneRegister RAM_OUT_101_F4_2_1   ( clk , write2_101  , RELUout_F4_2_1  , Final_101_F4_2_1  );
OneRegister RAM_OUT_101_F4_2_2   ( clk , write2_101  , RELUout_F4_2_2  , Final_101_F4_2_2  );
OneRegister RAM_OUT_102_F1_1_1   ( clk , write2_102  , RELUout_F1_1_1  , Final_102_F1_1_1  );
OneRegister RAM_OUT_102_F1_1_2   ( clk , write2_102  , RELUout_F1_1_2  , Final_102_F1_1_2  );
OneRegister RAM_OUT_102_F1_2_1   ( clk , write2_102  , RELUout_F1_2_1  , Final_102_F1_2_1  );
OneRegister RAM_OUT_102_F1_2_2   ( clk , write2_102  , RELUout_F1_2_2  , Final_102_F1_2_2  );
OneRegister RAM_OUT_102_F2_1_1   ( clk , write2_102  , RELUout_F2_1_1  , Final_102_F2_1_1  );
OneRegister RAM_OUT_102_F2_1_2   ( clk , write2_102  , RELUout_F2_1_2  , Final_102_F2_1_2  );
OneRegister RAM_OUT_102_F2_2_1   ( clk , write2_102  , RELUout_F2_2_1  , Final_102_F2_2_1  );
OneRegister RAM_OUT_102_F2_2_2   ( clk , write2_102  , RELUout_F2_2_2  , Final_102_F2_2_2  );
OneRegister RAM_OUT_102_F3_1_1   ( clk , write2_102  , RELUout_F3_1_1  , Final_102_F3_1_1  );
OneRegister RAM_OUT_102_F3_1_2   ( clk , write2_102  , RELUout_F3_1_2  , Final_102_F3_1_2  );
OneRegister RAM_OUT_102_F3_2_1   ( clk , write2_102  , RELUout_F3_2_1  , Final_102_F3_2_1  );
OneRegister RAM_OUT_102_F3_2_2   ( clk , write2_102  , RELUout_F3_2_2  , Final_102_F3_2_2  );
OneRegister RAM_OUT_102_F4_1_1   ( clk , write2_102  , RELUout_F4_1_1  , Final_102_F4_1_1  );
OneRegister RAM_OUT_102_F4_1_2   ( clk , write2_102  , RELUout_F4_1_2  , Final_102_F4_1_2  );
OneRegister RAM_OUT_102_F4_2_1   ( clk , write2_102  , RELUout_F4_2_1  , Final_102_F4_2_1  );
OneRegister RAM_OUT_102_F4_2_2   ( clk , write2_102  , RELUout_F4_2_2  , Final_102_F4_2_2  );
OneRegister RAM_OUT_103_F1_1_1   ( clk , write2_103  , RELUout_F1_1_1  , Final_103_F1_1_1  );
OneRegister RAM_OUT_103_F1_1_2   ( clk , write2_103  , RELUout_F1_1_2  , Final_103_F1_1_2  );
OneRegister RAM_OUT_103_F1_2_1   ( clk , write2_103  , RELUout_F1_2_1  , Final_103_F1_2_1  );
OneRegister RAM_OUT_103_F1_2_2   ( clk , write2_103  , RELUout_F1_2_2  , Final_103_F1_2_2  );
OneRegister RAM_OUT_103_F2_1_1   ( clk , write2_103  , RELUout_F2_1_1  , Final_103_F2_1_1  );
OneRegister RAM_OUT_103_F2_1_2   ( clk , write2_103  , RELUout_F2_1_2  , Final_103_F2_1_2  );
OneRegister RAM_OUT_103_F2_2_1   ( clk , write2_103  , RELUout_F2_2_1  , Final_103_F2_2_1  );
OneRegister RAM_OUT_103_F2_2_2   ( clk , write2_103  , RELUout_F2_2_2  , Final_103_F2_2_2  );
OneRegister RAM_OUT_103_F3_1_1   ( clk , write2_103  , RELUout_F3_1_1  , Final_103_F3_1_1  );
OneRegister RAM_OUT_103_F3_1_2   ( clk , write2_103  , RELUout_F3_1_2  , Final_103_F3_1_2  );
OneRegister RAM_OUT_103_F3_2_1   ( clk , write2_103  , RELUout_F3_2_1  , Final_103_F3_2_1  );
OneRegister RAM_OUT_103_F3_2_2   ( clk , write2_103  , RELUout_F3_2_2  , Final_103_F3_2_2  );
OneRegister RAM_OUT_103_F4_1_1   ( clk , write2_103  , RELUout_F4_1_1  , Final_103_F4_1_1  );
OneRegister RAM_OUT_103_F4_1_2   ( clk , write2_103  , RELUout_F4_1_2  , Final_103_F4_1_2  );
OneRegister RAM_OUT_103_F4_2_1   ( clk , write2_103  , RELUout_F4_2_1  , Final_103_F4_2_1  );
OneRegister RAM_OUT_103_F4_2_2   ( clk , write2_103  , RELUout_F4_2_2  , Final_103_F4_2_2  );
OneRegister RAM_OUT_104_F1_1_1   ( clk , write2_104  , RELUout_F1_1_1  , Final_104_F1_1_1  );
OneRegister RAM_OUT_104_F1_1_2   ( clk , write2_104  , RELUout_F1_1_2  , Final_104_F1_1_2  );
OneRegister RAM_OUT_104_F1_2_1   ( clk , write2_104  , RELUout_F1_2_1  , Final_104_F1_2_1  );
OneRegister RAM_OUT_104_F1_2_2   ( clk , write2_104  , RELUout_F1_2_2  , Final_104_F1_2_2  );
OneRegister RAM_OUT_104_F2_1_1   ( clk , write2_104  , RELUout_F2_1_1  , Final_104_F2_1_1  );
OneRegister RAM_OUT_104_F2_1_2   ( clk , write2_104  , RELUout_F2_1_2  , Final_104_F2_1_2  );
OneRegister RAM_OUT_104_F2_2_1   ( clk , write2_104  , RELUout_F2_2_1  , Final_104_F2_2_1  );
OneRegister RAM_OUT_104_F2_2_2   ( clk , write2_104  , RELUout_F2_2_2  , Final_104_F2_2_2  );
OneRegister RAM_OUT_104_F3_1_1   ( clk , write2_104  , RELUout_F3_1_1  , Final_104_F3_1_1  );
OneRegister RAM_OUT_104_F3_1_2   ( clk , write2_104  , RELUout_F3_1_2  , Final_104_F3_1_2  );
OneRegister RAM_OUT_104_F3_2_1   ( clk , write2_104  , RELUout_F3_2_1  , Final_104_F3_2_1  );
OneRegister RAM_OUT_104_F3_2_2   ( clk , write2_104  , RELUout_F3_2_2  , Final_104_F3_2_2  );
OneRegister RAM_OUT_104_F4_1_1   ( clk , write2_104  , RELUout_F4_1_1  , Final_104_F4_1_1  );
OneRegister RAM_OUT_104_F4_1_2   ( clk , write2_104  , RELUout_F4_1_2  , Final_104_F4_1_2  );
OneRegister RAM_OUT_104_F4_2_1   ( clk , write2_104  , RELUout_F4_2_1  , Final_104_F4_2_1  );
OneRegister RAM_OUT_104_F4_2_2   ( clk , write2_104  , RELUout_F4_2_2  , Final_104_F4_2_2  );
OneRegister RAM_OUT_105_F1_1_1   ( clk , write2_105  , RELUout_F1_1_1  , Final_105_F1_1_1  );
OneRegister RAM_OUT_105_F1_1_2   ( clk , write2_105  , RELUout_F1_1_2  , Final_105_F1_1_2  );
OneRegister RAM_OUT_105_F1_2_1   ( clk , write2_105  , RELUout_F1_2_1  , Final_105_F1_2_1  );
OneRegister RAM_OUT_105_F1_2_2   ( clk , write2_105  , RELUout_F1_2_2  , Final_105_F1_2_2  );
OneRegister RAM_OUT_105_F2_1_1   ( clk , write2_105  , RELUout_F2_1_1  , Final_105_F2_1_1  );
OneRegister RAM_OUT_105_F2_1_2   ( clk , write2_105  , RELUout_F2_1_2  , Final_105_F2_1_2  );
OneRegister RAM_OUT_105_F2_2_1   ( clk , write2_105  , RELUout_F2_2_1  , Final_105_F2_2_1  );
OneRegister RAM_OUT_105_F2_2_2   ( clk , write2_105  , RELUout_F2_2_2  , Final_105_F2_2_2  );
OneRegister RAM_OUT_105_F3_1_1   ( clk , write2_105  , RELUout_F3_1_1  , Final_105_F3_1_1  );
OneRegister RAM_OUT_105_F3_1_2   ( clk , write2_105  , RELUout_F3_1_2  , Final_105_F3_1_2  );
OneRegister RAM_OUT_105_F3_2_1   ( clk , write2_105  , RELUout_F3_2_1  , Final_105_F3_2_1  );
OneRegister RAM_OUT_105_F3_2_2   ( clk , write2_105  , RELUout_F3_2_2  , Final_105_F3_2_2  );
OneRegister RAM_OUT_105_F4_1_1   ( clk , write2_105  , RELUout_F4_1_1  , Final_105_F4_1_1  );
OneRegister RAM_OUT_105_F4_1_2   ( clk , write2_105  , RELUout_F4_1_2  , Final_105_F4_1_2  );
OneRegister RAM_OUT_105_F4_2_1   ( clk , write2_105  , RELUout_F4_2_1  , Final_105_F4_2_1  );
OneRegister RAM_OUT_105_F4_2_2   ( clk , write2_105  , RELUout_F4_2_2  , Final_105_F4_2_2  );
OneRegister RAM_OUT_106_F1_1_1   ( clk , write2_106  , RELUout_F1_1_1  , Final_106_F1_1_1  );
OneRegister RAM_OUT_106_F1_1_2   ( clk , write2_106  , RELUout_F1_1_2  , Final_106_F1_1_2  );
OneRegister RAM_OUT_106_F1_2_1   ( clk , write2_106  , RELUout_F1_2_1  , Final_106_F1_2_1  );
OneRegister RAM_OUT_106_F1_2_2   ( clk , write2_106  , RELUout_F1_2_2  , Final_106_F1_2_2  );
OneRegister RAM_OUT_106_F2_1_1   ( clk , write2_106  , RELUout_F2_1_1  , Final_106_F2_1_1  );
OneRegister RAM_OUT_106_F2_1_2   ( clk , write2_106  , RELUout_F2_1_2  , Final_106_F2_1_2  );
OneRegister RAM_OUT_106_F2_2_1   ( clk , write2_106  , RELUout_F2_2_1  , Final_106_F2_2_1  );
OneRegister RAM_OUT_106_F2_2_2   ( clk , write2_106  , RELUout_F2_2_2  , Final_106_F2_2_2  );
OneRegister RAM_OUT_106_F3_1_1   ( clk , write2_106  , RELUout_F3_1_1  , Final_106_F3_1_1  );
OneRegister RAM_OUT_106_F3_1_2   ( clk , write2_106  , RELUout_F3_1_2  , Final_106_F3_1_2  );
OneRegister RAM_OUT_106_F3_2_1   ( clk , write2_106  , RELUout_F3_2_1  , Final_106_F3_2_1  );
OneRegister RAM_OUT_106_F3_2_2   ( clk , write2_106  , RELUout_F3_2_2  , Final_106_F3_2_2  );
OneRegister RAM_OUT_106_F4_1_1   ( clk , write2_106  , RELUout_F4_1_1  , Final_106_F4_1_1  );
OneRegister RAM_OUT_106_F4_1_2   ( clk , write2_106  , RELUout_F4_1_2  , Final_106_F4_1_2  );
OneRegister RAM_OUT_106_F4_2_1   ( clk , write2_106  , RELUout_F4_2_1  , Final_106_F4_2_1  );
OneRegister RAM_OUT_106_F4_2_2   ( clk , write2_106  , RELUout_F4_2_2  , Final_106_F4_2_2  );
OneRegister RAM_OUT_107_F1_1_1   ( clk , write2_107  , RELUout_F1_1_1  , Final_107_F1_1_1  );
OneRegister RAM_OUT_107_F1_1_2   ( clk , write2_107  , RELUout_F1_1_2  , Final_107_F1_1_2  );
OneRegister RAM_OUT_107_F1_2_1   ( clk , write2_107  , RELUout_F1_2_1  , Final_107_F1_2_1  );
OneRegister RAM_OUT_107_F1_2_2   ( clk , write2_107  , RELUout_F1_2_2  , Final_107_F1_2_2  );
OneRegister RAM_OUT_107_F2_1_1   ( clk , write2_107  , RELUout_F2_1_1  , Final_107_F2_1_1  );
OneRegister RAM_OUT_107_F2_1_2   ( clk , write2_107  , RELUout_F2_1_2  , Final_107_F2_1_2  );
OneRegister RAM_OUT_107_F2_2_1   ( clk , write2_107  , RELUout_F2_2_1  , Final_107_F2_2_1  );
OneRegister RAM_OUT_107_F2_2_2   ( clk , write2_107  , RELUout_F2_2_2  , Final_107_F2_2_2  );
OneRegister RAM_OUT_107_F3_1_1   ( clk , write2_107  , RELUout_F3_1_1  , Final_107_F3_1_1  );
OneRegister RAM_OUT_107_F3_1_2   ( clk , write2_107  , RELUout_F3_1_2  , Final_107_F3_1_2  );
OneRegister RAM_OUT_107_F3_2_1   ( clk , write2_107  , RELUout_F3_2_1  , Final_107_F3_2_1  );
OneRegister RAM_OUT_107_F3_2_2   ( clk , write2_107  , RELUout_F3_2_2  , Final_107_F3_2_2  );
OneRegister RAM_OUT_107_F4_1_1   ( clk , write2_107  , RELUout_F4_1_1  , Final_107_F4_1_1  );
OneRegister RAM_OUT_107_F4_1_2   ( clk , write2_107  , RELUout_F4_1_2  , Final_107_F4_1_2  );
OneRegister RAM_OUT_107_F4_2_1   ( clk , write2_107  , RELUout_F4_2_1  , Final_107_F4_2_1  );
OneRegister RAM_OUT_107_F4_2_2   ( clk , write2_107  , RELUout_F4_2_2  , Final_107_F4_2_2  );
OneRegister RAM_OUT_108_F1_1_1   ( clk , write2_108  , RELUout_F1_1_1  , Final_108_F1_1_1  );
OneRegister RAM_OUT_108_F1_1_2   ( clk , write2_108  , RELUout_F1_1_2  , Final_108_F1_1_2  );
OneRegister RAM_OUT_108_F1_2_1   ( clk , write2_108  , RELUout_F1_2_1  , Final_108_F1_2_1  );
OneRegister RAM_OUT_108_F1_2_2   ( clk , write2_108  , RELUout_F1_2_2  , Final_108_F1_2_2  );
OneRegister RAM_OUT_108_F2_1_1   ( clk , write2_108  , RELUout_F2_1_1  , Final_108_F2_1_1  );
OneRegister RAM_OUT_108_F2_1_2   ( clk , write2_108  , RELUout_F2_1_2  , Final_108_F2_1_2  );
OneRegister RAM_OUT_108_F2_2_1   ( clk , write2_108  , RELUout_F2_2_1  , Final_108_F2_2_1  );
OneRegister RAM_OUT_108_F2_2_2   ( clk , write2_108  , RELUout_F2_2_2  , Final_108_F2_2_2  );
OneRegister RAM_OUT_108_F3_1_1   ( clk , write2_108  , RELUout_F3_1_1  , Final_108_F3_1_1  );
OneRegister RAM_OUT_108_F3_1_2   ( clk , write2_108  , RELUout_F3_1_2  , Final_108_F3_1_2  );
OneRegister RAM_OUT_108_F3_2_1   ( clk , write2_108  , RELUout_F3_2_1  , Final_108_F3_2_1  );
OneRegister RAM_OUT_108_F3_2_2   ( clk , write2_108  , RELUout_F3_2_2  , Final_108_F3_2_2  );
OneRegister RAM_OUT_108_F4_1_1   ( clk , write2_108  , RELUout_F4_1_1  , Final_108_F4_1_1  );
OneRegister RAM_OUT_108_F4_1_2   ( clk , write2_108  , RELUout_F4_1_2  , Final_108_F4_1_2  );
OneRegister RAM_OUT_108_F4_2_1   ( clk , write2_108  , RELUout_F4_2_1  , Final_108_F4_2_1  );
OneRegister RAM_OUT_108_F4_2_2   ( clk , write2_108  , RELUout_F4_2_2  , Final_108_F4_2_2  );
OneRegister RAM_OUT_109_F1_1_1   ( clk , write2_109  , RELUout_F1_1_1  , Final_109_F1_1_1  );
OneRegister RAM_OUT_109_F1_1_2   ( clk , write2_109  , RELUout_F1_1_2  , Final_109_F1_1_2  );
OneRegister RAM_OUT_109_F1_2_1   ( clk , write2_109  , RELUout_F1_2_1  , Final_109_F1_2_1  );
OneRegister RAM_OUT_109_F1_2_2   ( clk , write2_109  , RELUout_F1_2_2  , Final_109_F1_2_2  );
OneRegister RAM_OUT_109_F2_1_1   ( clk , write2_109  , RELUout_F2_1_1  , Final_109_F2_1_1  );
OneRegister RAM_OUT_109_F2_1_2   ( clk , write2_109  , RELUout_F2_1_2  , Final_109_F2_1_2  );
OneRegister RAM_OUT_109_F2_2_1   ( clk , write2_109  , RELUout_F2_2_1  , Final_109_F2_2_1  );
OneRegister RAM_OUT_109_F2_2_2   ( clk , write2_109  , RELUout_F2_2_2  , Final_109_F2_2_2  );
OneRegister RAM_OUT_109_F3_1_1   ( clk , write2_109  , RELUout_F3_1_1  , Final_109_F3_1_1  );
OneRegister RAM_OUT_109_F3_1_2   ( clk , write2_109  , RELUout_F3_1_2  , Final_109_F3_1_2  );
OneRegister RAM_OUT_109_F3_2_1   ( clk , write2_109  , RELUout_F3_2_1  , Final_109_F3_2_1  );
OneRegister RAM_OUT_109_F3_2_2   ( clk , write2_109  , RELUout_F3_2_2  , Final_109_F3_2_2  );
OneRegister RAM_OUT_109_F4_1_1   ( clk , write2_109  , RELUout_F4_1_1  , Final_109_F4_1_1  );
OneRegister RAM_OUT_109_F4_1_2   ( clk , write2_109  , RELUout_F4_1_2  , Final_109_F4_1_2  );
OneRegister RAM_OUT_109_F4_2_1   ( clk , write2_109  , RELUout_F4_2_1  , Final_109_F4_2_1  );
OneRegister RAM_OUT_109_F4_2_2   ( clk , write2_109  , RELUout_F4_2_2  , Final_109_F4_2_2  );
OneRegister RAM_OUT_110_F1_1_1   ( clk , write2_110  , RELUout_F1_1_1  , Final_110_F1_1_1  );
OneRegister RAM_OUT_110_F1_1_2   ( clk , write2_110  , RELUout_F1_1_2  , Final_110_F1_1_2  );
OneRegister RAM_OUT_110_F1_2_1   ( clk , write2_110  , RELUout_F1_2_1  , Final_110_F1_2_1  );
OneRegister RAM_OUT_110_F1_2_2   ( clk , write2_110  , RELUout_F1_2_2  , Final_110_F1_2_2  );
OneRegister RAM_OUT_110_F2_1_1   ( clk , write2_110  , RELUout_F2_1_1  , Final_110_F2_1_1  );
OneRegister RAM_OUT_110_F2_1_2   ( clk , write2_110  , RELUout_F2_1_2  , Final_110_F2_1_2  );
OneRegister RAM_OUT_110_F2_2_1   ( clk , write2_110  , RELUout_F2_2_1  , Final_110_F2_2_1  );
OneRegister RAM_OUT_110_F2_2_2   ( clk , write2_110  , RELUout_F2_2_2  , Final_110_F2_2_2  );
OneRegister RAM_OUT_110_F3_1_1   ( clk , write2_110  , RELUout_F3_1_1  , Final_110_F3_1_1  );
OneRegister RAM_OUT_110_F3_1_2   ( clk , write2_110  , RELUout_F3_1_2  , Final_110_F3_1_2  );
OneRegister RAM_OUT_110_F3_2_1   ( clk , write2_110  , RELUout_F3_2_1  , Final_110_F3_2_1  );
OneRegister RAM_OUT_110_F3_2_2   ( clk , write2_110  , RELUout_F3_2_2  , Final_110_F3_2_2  );
OneRegister RAM_OUT_110_F4_1_1   ( clk , write2_110  , RELUout_F4_1_1  , Final_110_F4_1_1  );
OneRegister RAM_OUT_110_F4_1_2   ( clk , write2_110  , RELUout_F4_1_2  , Final_110_F4_1_2  );
OneRegister RAM_OUT_110_F4_2_1   ( clk , write2_110  , RELUout_F4_2_1  , Final_110_F4_2_1  );
OneRegister RAM_OUT_110_F4_2_2   ( clk , write2_110  , RELUout_F4_2_2  , Final_110_F4_2_2  );
OneRegister RAM_OUT_111_F1_1_1   ( clk , write2_111  , RELUout_F1_1_1  , Final_111_F1_1_1  );
OneRegister RAM_OUT_111_F1_1_2   ( clk , write2_111  , RELUout_F1_1_2  , Final_111_F1_1_2  );
OneRegister RAM_OUT_111_F1_2_1   ( clk , write2_111  , RELUout_F1_2_1  , Final_111_F1_2_1  );
OneRegister RAM_OUT_111_F1_2_2   ( clk , write2_111  , RELUout_F1_2_2  , Final_111_F1_2_2  );
OneRegister RAM_OUT_111_F2_1_1   ( clk , write2_111  , RELUout_F2_1_1  , Final_111_F2_1_1  );
OneRegister RAM_OUT_111_F2_1_2   ( clk , write2_111  , RELUout_F2_1_2  , Final_111_F2_1_2  );
OneRegister RAM_OUT_111_F2_2_1   ( clk , write2_111  , RELUout_F2_2_1  , Final_111_F2_2_1  );
OneRegister RAM_OUT_111_F2_2_2   ( clk , write2_111  , RELUout_F2_2_2  , Final_111_F2_2_2  );
OneRegister RAM_OUT_111_F3_1_1   ( clk , write2_111  , RELUout_F3_1_1  , Final_111_F3_1_1  );
OneRegister RAM_OUT_111_F3_1_2   ( clk , write2_111  , RELUout_F3_1_2  , Final_111_F3_1_2  );
OneRegister RAM_OUT_111_F3_2_1   ( clk , write2_111  , RELUout_F3_2_1  , Final_111_F3_2_1  );
OneRegister RAM_OUT_111_F3_2_2   ( clk , write2_111  , RELUout_F3_2_2  , Final_111_F3_2_2  );
OneRegister RAM_OUT_111_F4_1_1   ( clk , write2_111  , RELUout_F4_1_1  , Final_111_F4_1_1  );
OneRegister RAM_OUT_111_F4_1_2   ( clk , write2_111  , RELUout_F4_1_2  , Final_111_F4_1_2  );
OneRegister RAM_OUT_111_F4_2_1   ( clk , write2_111  , RELUout_F4_2_1  , Final_111_F4_2_1  );
OneRegister RAM_OUT_111_F4_2_2   ( clk , write2_111  , RELUout_F4_2_2  , Final_111_F4_2_2  );
OneRegister RAM_OUT_112_F1_1_1   ( clk , write2_112  , RELUout_F1_1_1  , Final_112_F1_1_1  );
OneRegister RAM_OUT_112_F1_1_2   ( clk , write2_112  , RELUout_F1_1_2  , Final_112_F1_1_2  );
OneRegister RAM_OUT_112_F1_2_1   ( clk , write2_112  , RELUout_F1_2_1  , Final_112_F1_2_1  );
OneRegister RAM_OUT_112_F1_2_2   ( clk , write2_112  , RELUout_F1_2_2  , Final_112_F1_2_2  );
OneRegister RAM_OUT_112_F2_1_1   ( clk , write2_112  , RELUout_F2_1_1  , Final_112_F2_1_1  );
OneRegister RAM_OUT_112_F2_1_2   ( clk , write2_112  , RELUout_F2_1_2  , Final_112_F2_1_2  );
OneRegister RAM_OUT_112_F2_2_1   ( clk , write2_112  , RELUout_F2_2_1  , Final_112_F2_2_1  );
OneRegister RAM_OUT_112_F2_2_2   ( clk , write2_112  , RELUout_F2_2_2  , Final_112_F2_2_2  );
OneRegister RAM_OUT_112_F3_1_1   ( clk , write2_112  , RELUout_F3_1_1  , Final_112_F3_1_1  );
OneRegister RAM_OUT_112_F3_1_2   ( clk , write2_112  , RELUout_F3_1_2  , Final_112_F3_1_2  );
OneRegister RAM_OUT_112_F3_2_1   ( clk , write2_112  , RELUout_F3_2_1  , Final_112_F3_2_1  );
OneRegister RAM_OUT_112_F3_2_2   ( clk , write2_112  , RELUout_F3_2_2  , Final_112_F3_2_2  );
OneRegister RAM_OUT_112_F4_1_1   ( clk , write2_112  , RELUout_F4_1_1  , Final_112_F4_1_1  );
OneRegister RAM_OUT_112_F4_1_2   ( clk , write2_112  , RELUout_F4_1_2  , Final_112_F4_1_2  );
OneRegister RAM_OUT_112_F4_2_1   ( clk , write2_112  , RELUout_F4_2_1  , Final_112_F4_2_1  );
OneRegister RAM_OUT_112_F4_2_2   ( clk , write2_112  , RELUout_F4_2_2  , Final_112_F4_2_2  );
OneRegister RAM_OUT_113_F1_1_1   ( clk , write2_113  , RELUout_F1_1_1  , Final_113_F1_1_1  );
OneRegister RAM_OUT_113_F1_1_2   ( clk , write2_113  , RELUout_F1_1_2  , Final_113_F1_1_2  );
OneRegister RAM_OUT_113_F1_2_1   ( clk , write2_113  , RELUout_F1_2_1  , Final_113_F1_2_1  );
OneRegister RAM_OUT_113_F1_2_2   ( clk , write2_113  , RELUout_F1_2_2  , Final_113_F1_2_2  );
OneRegister RAM_OUT_113_F2_1_1   ( clk , write2_113  , RELUout_F2_1_1  , Final_113_F2_1_1  );
OneRegister RAM_OUT_113_F2_1_2   ( clk , write2_113  , RELUout_F2_1_2  , Final_113_F2_1_2  );
OneRegister RAM_OUT_113_F2_2_1   ( clk , write2_113  , RELUout_F2_2_1  , Final_113_F2_2_1  );
OneRegister RAM_OUT_113_F2_2_2   ( clk , write2_113  , RELUout_F2_2_2  , Final_113_F2_2_2  );
OneRegister RAM_OUT_113_F3_1_1   ( clk , write2_113  , RELUout_F3_1_1  , Final_113_F3_1_1  );
OneRegister RAM_OUT_113_F3_1_2   ( clk , write2_113  , RELUout_F3_1_2  , Final_113_F3_1_2  );
OneRegister RAM_OUT_113_F3_2_1   ( clk , write2_113  , RELUout_F3_2_1  , Final_113_F3_2_1  );
OneRegister RAM_OUT_113_F3_2_2   ( clk , write2_113  , RELUout_F3_2_2  , Final_113_F3_2_2  );
OneRegister RAM_OUT_113_F4_1_1   ( clk , write2_113  , RELUout_F4_1_1  , Final_113_F4_1_1  );
OneRegister RAM_OUT_113_F4_1_2   ( clk , write2_113  , RELUout_F4_1_2  , Final_113_F4_1_2  );
OneRegister RAM_OUT_113_F4_2_1   ( clk , write2_113  , RELUout_F4_2_1  , Final_113_F4_2_1  );
OneRegister RAM_OUT_113_F4_2_2   ( clk , write2_113  , RELUout_F4_2_2  , Final_113_F4_2_2  );
OneRegister RAM_OUT_114_F1_1_1   ( clk , write2_114  , RELUout_F1_1_1  , Final_114_F1_1_1  );
OneRegister RAM_OUT_114_F1_1_2   ( clk , write2_114  , RELUout_F1_1_2  , Final_114_F1_1_2  );
OneRegister RAM_OUT_114_F1_2_1   ( clk , write2_114  , RELUout_F1_2_1  , Final_114_F1_2_1  );
OneRegister RAM_OUT_114_F1_2_2   ( clk , write2_114  , RELUout_F1_2_2  , Final_114_F1_2_2  );
OneRegister RAM_OUT_114_F2_1_1   ( clk , write2_114  , RELUout_F2_1_1  , Final_114_F2_1_1  );
OneRegister RAM_OUT_114_F2_1_2   ( clk , write2_114  , RELUout_F2_1_2  , Final_114_F2_1_2  );
OneRegister RAM_OUT_114_F2_2_1   ( clk , write2_114  , RELUout_F2_2_1  , Final_114_F2_2_1  );
OneRegister RAM_OUT_114_F2_2_2   ( clk , write2_114  , RELUout_F2_2_2  , Final_114_F2_2_2  );
OneRegister RAM_OUT_114_F3_1_1   ( clk , write2_114  , RELUout_F3_1_1  , Final_114_F3_1_1  );
OneRegister RAM_OUT_114_F3_1_2   ( clk , write2_114  , RELUout_F3_1_2  , Final_114_F3_1_2  );
OneRegister RAM_OUT_114_F3_2_1   ( clk , write2_114  , RELUout_F3_2_1  , Final_114_F3_2_1  );
OneRegister RAM_OUT_114_F3_2_2   ( clk , write2_114  , RELUout_F3_2_2  , Final_114_F3_2_2  );
OneRegister RAM_OUT_114_F4_1_1   ( clk , write2_114  , RELUout_F4_1_1  , Final_114_F4_1_1  );
OneRegister RAM_OUT_114_F4_1_2   ( clk , write2_114  , RELUout_F4_1_2  , Final_114_F4_1_2  );
OneRegister RAM_OUT_114_F4_2_1   ( clk , write2_114  , RELUout_F4_2_1  , Final_114_F4_2_1  );
OneRegister RAM_OUT_114_F4_2_2   ( clk , write2_114  , RELUout_F4_2_2  , Final_114_F4_2_2  );
OneRegister RAM_OUT_115_F1_1_1   ( clk , write2_115  , RELUout_F1_1_1  , Final_115_F1_1_1  );
OneRegister RAM_OUT_115_F1_1_2   ( clk , write2_115  , RELUout_F1_1_2  , Final_115_F1_1_2  );
OneRegister RAM_OUT_115_F1_2_1   ( clk , write2_115  , RELUout_F1_2_1  , Final_115_F1_2_1  );
OneRegister RAM_OUT_115_F1_2_2   ( clk , write2_115  , RELUout_F1_2_2  , Final_115_F1_2_2  );
OneRegister RAM_OUT_115_F2_1_1   ( clk , write2_115  , RELUout_F2_1_1  , Final_115_F2_1_1  );
OneRegister RAM_OUT_115_F2_1_2   ( clk , write2_115  , RELUout_F2_1_2  , Final_115_F2_1_2  );
OneRegister RAM_OUT_115_F2_2_1   ( clk , write2_115  , RELUout_F2_2_1  , Final_115_F2_2_1  );
OneRegister RAM_OUT_115_F2_2_2   ( clk , write2_115  , RELUout_F2_2_2  , Final_115_F2_2_2  );
OneRegister RAM_OUT_115_F3_1_1   ( clk , write2_115  , RELUout_F3_1_1  , Final_115_F3_1_1  );
OneRegister RAM_OUT_115_F3_1_2   ( clk , write2_115  , RELUout_F3_1_2  , Final_115_F3_1_2  );
OneRegister RAM_OUT_115_F3_2_1   ( clk , write2_115  , RELUout_F3_2_1  , Final_115_F3_2_1  );
OneRegister RAM_OUT_115_F3_2_2   ( clk , write2_115  , RELUout_F3_2_2  , Final_115_F3_2_2  );
OneRegister RAM_OUT_115_F4_1_1   ( clk , write2_115  , RELUout_F4_1_1  , Final_115_F4_1_1  );
OneRegister RAM_OUT_115_F4_1_2   ( clk , write2_115  , RELUout_F4_1_2  , Final_115_F4_1_2  );
OneRegister RAM_OUT_115_F4_2_1   ( clk , write2_115  , RELUout_F4_2_1  , Final_115_F4_2_1  );
OneRegister RAM_OUT_115_F4_2_2   ( clk , write2_115  , RELUout_F4_2_2  , Final_115_F4_2_2  );
OneRegister RAM_OUT_116_F1_1_1   ( clk , write2_116  , RELUout_F1_1_1  , Final_116_F1_1_1  );
OneRegister RAM_OUT_116_F1_1_2   ( clk , write2_116  , RELUout_F1_1_2  , Final_116_F1_1_2  );
OneRegister RAM_OUT_116_F1_2_1   ( clk , write2_116  , RELUout_F1_2_1  , Final_116_F1_2_1  );
OneRegister RAM_OUT_116_F1_2_2   ( clk , write2_116  , RELUout_F1_2_2  , Final_116_F1_2_2  );
OneRegister RAM_OUT_116_F2_1_1   ( clk , write2_116  , RELUout_F2_1_1  , Final_116_F2_1_1  );
OneRegister RAM_OUT_116_F2_1_2   ( clk , write2_116  , RELUout_F2_1_2  , Final_116_F2_1_2  );
OneRegister RAM_OUT_116_F2_2_1   ( clk , write2_116  , RELUout_F2_2_1  , Final_116_F2_2_1  );
OneRegister RAM_OUT_116_F2_2_2   ( clk , write2_116  , RELUout_F2_2_2  , Final_116_F2_2_2  );
OneRegister RAM_OUT_116_F3_1_1   ( clk , write2_116  , RELUout_F3_1_1  , Final_116_F3_1_1  );
OneRegister RAM_OUT_116_F3_1_2   ( clk , write2_116  , RELUout_F3_1_2  , Final_116_F3_1_2  );
OneRegister RAM_OUT_116_F3_2_1   ( clk , write2_116  , RELUout_F3_2_1  , Final_116_F3_2_1  );
OneRegister RAM_OUT_116_F3_2_2   ( clk , write2_116  , RELUout_F3_2_2  , Final_116_F3_2_2  );
OneRegister RAM_OUT_116_F4_1_1   ( clk , write2_116  , RELUout_F4_1_1  , Final_116_F4_1_1  );
OneRegister RAM_OUT_116_F4_1_2   ( clk , write2_116  , RELUout_F4_1_2  , Final_116_F4_1_2  );
OneRegister RAM_OUT_116_F4_2_1   ( clk , write2_116  , RELUout_F4_2_1  , Final_116_F4_2_1  );
OneRegister RAM_OUT_116_F4_2_2   ( clk , write2_116  , RELUout_F4_2_2  , Final_116_F4_2_2  );
OneRegister RAM_OUT_117_F1_1_1   ( clk , write2_117  , RELUout_F1_1_1  , Final_117_F1_1_1  );
OneRegister RAM_OUT_117_F1_1_2   ( clk , write2_117  , RELUout_F1_1_2  , Final_117_F1_1_2  );
OneRegister RAM_OUT_117_F1_2_1   ( clk , write2_117  , RELUout_F1_2_1  , Final_117_F1_2_1  );
OneRegister RAM_OUT_117_F1_2_2   ( clk , write2_117  , RELUout_F1_2_2  , Final_117_F1_2_2  );
OneRegister RAM_OUT_117_F2_1_1   ( clk , write2_117  , RELUout_F2_1_1  , Final_117_F2_1_1  );
OneRegister RAM_OUT_117_F2_1_2   ( clk , write2_117  , RELUout_F2_1_2  , Final_117_F2_1_2  );
OneRegister RAM_OUT_117_F2_2_1   ( clk , write2_117  , RELUout_F2_2_1  , Final_117_F2_2_1  );
OneRegister RAM_OUT_117_F2_2_2   ( clk , write2_117  , RELUout_F2_2_2  , Final_117_F2_2_2  );
OneRegister RAM_OUT_117_F3_1_1   ( clk , write2_117  , RELUout_F3_1_1  , Final_117_F3_1_1  );
OneRegister RAM_OUT_117_F3_1_2   ( clk , write2_117  , RELUout_F3_1_2  , Final_117_F3_1_2  );
OneRegister RAM_OUT_117_F3_2_1   ( clk , write2_117  , RELUout_F3_2_1  , Final_117_F3_2_1  );
OneRegister RAM_OUT_117_F3_2_2   ( clk , write2_117  , RELUout_F3_2_2  , Final_117_F3_2_2  );
OneRegister RAM_OUT_117_F4_1_1   ( clk , write2_117  , RELUout_F4_1_1  , Final_117_F4_1_1  );
OneRegister RAM_OUT_117_F4_1_2   ( clk , write2_117  , RELUout_F4_1_2  , Final_117_F4_1_2  );
OneRegister RAM_OUT_117_F4_2_1   ( clk , write2_117  , RELUout_F4_2_1  , Final_117_F4_2_1  );
OneRegister RAM_OUT_117_F4_2_2   ( clk , write2_117  , RELUout_F4_2_2  , Final_117_F4_2_2  );
OneRegister RAM_OUT_118_F1_1_1   ( clk , write2_118  , RELUout_F1_1_1  , Final_118_F1_1_1  );
OneRegister RAM_OUT_118_F1_1_2   ( clk , write2_118  , RELUout_F1_1_2  , Final_118_F1_1_2  );
OneRegister RAM_OUT_118_F1_2_1   ( clk , write2_118  , RELUout_F1_2_1  , Final_118_F1_2_1  );
OneRegister RAM_OUT_118_F1_2_2   ( clk , write2_118  , RELUout_F1_2_2  , Final_118_F1_2_2  );
OneRegister RAM_OUT_118_F2_1_1   ( clk , write2_118  , RELUout_F2_1_1  , Final_118_F2_1_1  );
OneRegister RAM_OUT_118_F2_1_2   ( clk , write2_118  , RELUout_F2_1_2  , Final_118_F2_1_2  );
OneRegister RAM_OUT_118_F2_2_1   ( clk , write2_118  , RELUout_F2_2_1  , Final_118_F2_2_1  );
OneRegister RAM_OUT_118_F2_2_2   ( clk , write2_118  , RELUout_F2_2_2  , Final_118_F2_2_2  );
OneRegister RAM_OUT_118_F3_1_1   ( clk , write2_118  , RELUout_F3_1_1  , Final_118_F3_1_1  );
OneRegister RAM_OUT_118_F3_1_2   ( clk , write2_118  , RELUout_F3_1_2  , Final_118_F3_1_2  );
OneRegister RAM_OUT_118_F3_2_1   ( clk , write2_118  , RELUout_F3_2_1  , Final_118_F3_2_1  );
OneRegister RAM_OUT_118_F3_2_2   ( clk , write2_118  , RELUout_F3_2_2  , Final_118_F3_2_2  );
OneRegister RAM_OUT_118_F4_1_1   ( clk , write2_118  , RELUout_F4_1_1  , Final_118_F4_1_1  );
OneRegister RAM_OUT_118_F4_1_2   ( clk , write2_118  , RELUout_F4_1_2  , Final_118_F4_1_2  );
OneRegister RAM_OUT_118_F4_2_1   ( clk , write2_118  , RELUout_F4_2_1  , Final_118_F4_2_1  );
OneRegister RAM_OUT_118_F4_2_2   ( clk , write2_118  , RELUout_F4_2_2  , Final_118_F4_2_2  );
OneRegister RAM_OUT_119_F1_1_1   ( clk , write2_119  , RELUout_F1_1_1  , Final_119_F1_1_1  );
OneRegister RAM_OUT_119_F1_1_2   ( clk , write2_119  , RELUout_F1_1_2  , Final_119_F1_1_2  );
OneRegister RAM_OUT_119_F1_2_1   ( clk , write2_119  , RELUout_F1_2_1  , Final_119_F1_2_1  );
OneRegister RAM_OUT_119_F1_2_2   ( clk , write2_119  , RELUout_F1_2_2  , Final_119_F1_2_2  );
OneRegister RAM_OUT_119_F2_1_1   ( clk , write2_119  , RELUout_F2_1_1  , Final_119_F2_1_1  );
OneRegister RAM_OUT_119_F2_1_2   ( clk , write2_119  , RELUout_F2_1_2  , Final_119_F2_1_2  );
OneRegister RAM_OUT_119_F2_2_1   ( clk , write2_119  , RELUout_F2_2_1  , Final_119_F2_2_1  );
OneRegister RAM_OUT_119_F2_2_2   ( clk , write2_119  , RELUout_F2_2_2  , Final_119_F2_2_2  );
OneRegister RAM_OUT_119_F3_1_1   ( clk , write2_119  , RELUout_F3_1_1  , Final_119_F3_1_1  );
OneRegister RAM_OUT_119_F3_1_2   ( clk , write2_119  , RELUout_F3_1_2  , Final_119_F3_1_2  );
OneRegister RAM_OUT_119_F3_2_1   ( clk , write2_119  , RELUout_F3_2_1  , Final_119_F3_2_1  );
OneRegister RAM_OUT_119_F3_2_2   ( clk , write2_119  , RELUout_F3_2_2  , Final_119_F3_2_2  );
OneRegister RAM_OUT_119_F4_1_1   ( clk , write2_119  , RELUout_F4_1_1  , Final_119_F4_1_1  );
OneRegister RAM_OUT_119_F4_1_2   ( clk , write2_119  , RELUout_F4_1_2  , Final_119_F4_1_2  );
OneRegister RAM_OUT_119_F4_2_1   ( clk , write2_119  , RELUout_F4_2_1  , Final_119_F4_2_1  );
OneRegister RAM_OUT_119_F4_2_2   ( clk , write2_119  , RELUout_F4_2_2  , Final_119_F4_2_2  );
OneRegister RAM_OUT_120_F1_1_1   ( clk , write2_120  , RELUout_F1_1_1  , Final_120_F1_1_1  );
OneRegister RAM_OUT_120_F1_1_2   ( clk , write2_120  , RELUout_F1_1_2  , Final_120_F1_1_2  );
OneRegister RAM_OUT_120_F1_2_1   ( clk , write2_120  , RELUout_F1_2_1  , Final_120_F1_2_1  );
OneRegister RAM_OUT_120_F1_2_2   ( clk , write2_120  , RELUout_F1_2_2  , Final_120_F1_2_2  );
OneRegister RAM_OUT_120_F2_1_1   ( clk , write2_120  , RELUout_F2_1_1  , Final_120_F2_1_1  );
OneRegister RAM_OUT_120_F2_1_2   ( clk , write2_120  , RELUout_F2_1_2  , Final_120_F2_1_2  );
OneRegister RAM_OUT_120_F2_2_1   ( clk , write2_120  , RELUout_F2_2_1  , Final_120_F2_2_1  );
OneRegister RAM_OUT_120_F2_2_2   ( clk , write2_120  , RELUout_F2_2_2  , Final_120_F2_2_2  );
OneRegister RAM_OUT_120_F3_1_1   ( clk , write2_120  , RELUout_F3_1_1  , Final_120_F3_1_1  );
OneRegister RAM_OUT_120_F3_1_2   ( clk , write2_120  , RELUout_F3_1_2  , Final_120_F3_1_2  );
OneRegister RAM_OUT_120_F3_2_1   ( clk , write2_120  , RELUout_F3_2_1  , Final_120_F3_2_1  );
OneRegister RAM_OUT_120_F3_2_2   ( clk , write2_120  , RELUout_F3_2_2  , Final_120_F3_2_2  );
OneRegister RAM_OUT_120_F4_1_1   ( clk , write2_120  , RELUout_F4_1_1  , Final_120_F4_1_1  );
OneRegister RAM_OUT_120_F4_1_2   ( clk , write2_120  , RELUout_F4_1_2  , Final_120_F4_1_2  );
OneRegister RAM_OUT_120_F4_2_1   ( clk , write2_120  , RELUout_F4_2_1  , Final_120_F4_2_1  );
OneRegister RAM_OUT_120_F4_2_2   ( clk , write2_120  , RELUout_F4_2_2  , Final_120_F4_2_2  );
OneRegister RAM_OUT_121_F1_1_1   ( clk , write2_121  , RELUout_F1_1_1  , Final_121_F1_1_1  );
OneRegister RAM_OUT_121_F1_1_2   ( clk , write2_121  , RELUout_F1_1_2  , Final_121_F1_1_2  );
OneRegister RAM_OUT_121_F1_2_1   ( clk , write2_121  , RELUout_F1_2_1  , Final_121_F1_2_1  );
OneRegister RAM_OUT_121_F1_2_2   ( clk , write2_121  , RELUout_F1_2_2  , Final_121_F1_2_2  );
OneRegister RAM_OUT_121_F2_1_1   ( clk , write2_121  , RELUout_F2_1_1  , Final_121_F2_1_1  );
OneRegister RAM_OUT_121_F2_1_2   ( clk , write2_121  , RELUout_F2_1_2  , Final_121_F2_1_2  );
OneRegister RAM_OUT_121_F2_2_1   ( clk , write2_121  , RELUout_F2_2_1  , Final_121_F2_2_1  );
OneRegister RAM_OUT_121_F2_2_2   ( clk , write2_121  , RELUout_F2_2_2  , Final_121_F2_2_2  );
OneRegister RAM_OUT_121_F3_1_1   ( clk , write2_121  , RELUout_F3_1_1  , Final_121_F3_1_1  );
OneRegister RAM_OUT_121_F3_1_2   ( clk , write2_121  , RELUout_F3_1_2  , Final_121_F3_1_2  );
OneRegister RAM_OUT_121_F3_2_1   ( clk , write2_121  , RELUout_F3_2_1  , Final_121_F3_2_1  );
OneRegister RAM_OUT_121_F3_2_2   ( clk , write2_121  , RELUout_F3_2_2  , Final_121_F3_2_2  );
OneRegister RAM_OUT_121_F4_1_1   ( clk , write2_121  , RELUout_F4_1_1  , Final_121_F4_1_1  );
OneRegister RAM_OUT_121_F4_1_2   ( clk , write2_121  , RELUout_F4_1_2  , Final_121_F4_1_2  );
OneRegister RAM_OUT_121_F4_2_1   ( clk , write2_121  , RELUout_F4_2_1  , Final_121_F4_2_1  );
OneRegister RAM_OUT_121_F4_2_2   ( clk , write2_121  , RELUout_F4_2_2  , Final_121_F4_2_2  );
OneRegister RAM_OUT_122_F1_1_1   ( clk , write2_122  , RELUout_F1_1_1  , Final_122_F1_1_1  );
OneRegister RAM_OUT_122_F1_1_2   ( clk , write2_122  , RELUout_F1_1_2  , Final_122_F1_1_2  );
OneRegister RAM_OUT_122_F1_2_1   ( clk , write2_122  , RELUout_F1_2_1  , Final_122_F1_2_1  );
OneRegister RAM_OUT_122_F1_2_2   ( clk , write2_122  , RELUout_F1_2_2  , Final_122_F1_2_2  );
OneRegister RAM_OUT_122_F2_1_1   ( clk , write2_122  , RELUout_F2_1_1  , Final_122_F2_1_1  );
OneRegister RAM_OUT_122_F2_1_2   ( clk , write2_122  , RELUout_F2_1_2  , Final_122_F2_1_2  );
OneRegister RAM_OUT_122_F2_2_1   ( clk , write2_122  , RELUout_F2_2_1  , Final_122_F2_2_1  );
OneRegister RAM_OUT_122_F2_2_2   ( clk , write2_122  , RELUout_F2_2_2  , Final_122_F2_2_2  );
OneRegister RAM_OUT_122_F3_1_1   ( clk , write2_122  , RELUout_F3_1_1  , Final_122_F3_1_1  );
OneRegister RAM_OUT_122_F3_1_2   ( clk , write2_122  , RELUout_F3_1_2  , Final_122_F3_1_2  );
OneRegister RAM_OUT_122_F3_2_1   ( clk , write2_122  , RELUout_F3_2_1  , Final_122_F3_2_1  );
OneRegister RAM_OUT_122_F3_2_2   ( clk , write2_122  , RELUout_F3_2_2  , Final_122_F3_2_2  );
OneRegister RAM_OUT_122_F4_1_1   ( clk , write2_122  , RELUout_F4_1_1  , Final_122_F4_1_1  );
OneRegister RAM_OUT_122_F4_1_2   ( clk , write2_122  , RELUout_F4_1_2  , Final_122_F4_1_2  );
OneRegister RAM_OUT_122_F4_2_1   ( clk , write2_122  , RELUout_F4_2_1  , Final_122_F4_2_1  );
OneRegister RAM_OUT_122_F4_2_2   ( clk , write2_122  , RELUout_F4_2_2  , Final_122_F4_2_2  );
OneRegister RAM_OUT_123_F1_1_1   ( clk , write2_123  , RELUout_F1_1_1  , Final_123_F1_1_1  );
OneRegister RAM_OUT_123_F1_1_2   ( clk , write2_123  , RELUout_F1_1_2  , Final_123_F1_1_2  );
OneRegister RAM_OUT_123_F1_2_1   ( clk , write2_123  , RELUout_F1_2_1  , Final_123_F1_2_1  );
OneRegister RAM_OUT_123_F1_2_2   ( clk , write2_123  , RELUout_F1_2_2  , Final_123_F1_2_2  );
OneRegister RAM_OUT_123_F2_1_1   ( clk , write2_123  , RELUout_F2_1_1  , Final_123_F2_1_1  );
OneRegister RAM_OUT_123_F2_1_2   ( clk , write2_123  , RELUout_F2_1_2  , Final_123_F2_1_2  );
OneRegister RAM_OUT_123_F2_2_1   ( clk , write2_123  , RELUout_F2_2_1  , Final_123_F2_2_1  );
OneRegister RAM_OUT_123_F2_2_2   ( clk , write2_123  , RELUout_F2_2_2  , Final_123_F2_2_2  );
OneRegister RAM_OUT_123_F3_1_1   ( clk , write2_123  , RELUout_F3_1_1  , Final_123_F3_1_1  );
OneRegister RAM_OUT_123_F3_1_2   ( clk , write2_123  , RELUout_F3_1_2  , Final_123_F3_1_2  );
OneRegister RAM_OUT_123_F3_2_1   ( clk , write2_123  , RELUout_F3_2_1  , Final_123_F3_2_1  );
OneRegister RAM_OUT_123_F3_2_2   ( clk , write2_123  , RELUout_F3_2_2  , Final_123_F3_2_2  );
OneRegister RAM_OUT_123_F4_1_1   ( clk , write2_123  , RELUout_F4_1_1  , Final_123_F4_1_1  );
OneRegister RAM_OUT_123_F4_1_2   ( clk , write2_123  , RELUout_F4_1_2  , Final_123_F4_1_2  );
OneRegister RAM_OUT_123_F4_2_1   ( clk , write2_123  , RELUout_F4_2_1  , Final_123_F4_2_1  );
OneRegister RAM_OUT_123_F4_2_2   ( clk , write2_123  , RELUout_F4_2_2  , Final_123_F4_2_2  );
OneRegister RAM_OUT_124_F1_1_1   ( clk , write2_124  , RELUout_F1_1_1  , Final_124_F1_1_1  );
OneRegister RAM_OUT_124_F1_1_2   ( clk , write2_124  , RELUout_F1_1_2  , Final_124_F1_1_2  );
OneRegister RAM_OUT_124_F1_2_1   ( clk , write2_124  , RELUout_F1_2_1  , Final_124_F1_2_1  );
OneRegister RAM_OUT_124_F1_2_2   ( clk , write2_124  , RELUout_F1_2_2  , Final_124_F1_2_2  );
OneRegister RAM_OUT_124_F2_1_1   ( clk , write2_124  , RELUout_F2_1_1  , Final_124_F2_1_1  );
OneRegister RAM_OUT_124_F2_1_2   ( clk , write2_124  , RELUout_F2_1_2  , Final_124_F2_1_2  );
OneRegister RAM_OUT_124_F2_2_1   ( clk , write2_124  , RELUout_F2_2_1  , Final_124_F2_2_1  );
OneRegister RAM_OUT_124_F2_2_2   ( clk , write2_124  , RELUout_F2_2_2  , Final_124_F2_2_2  );
OneRegister RAM_OUT_124_F3_1_1   ( clk , write2_124  , RELUout_F3_1_1  , Final_124_F3_1_1  );
OneRegister RAM_OUT_124_F3_1_2   ( clk , write2_124  , RELUout_F3_1_2  , Final_124_F3_1_2  );
OneRegister RAM_OUT_124_F3_2_1   ( clk , write2_124  , RELUout_F3_2_1  , Final_124_F3_2_1  );
OneRegister RAM_OUT_124_F3_2_2   ( clk , write2_124  , RELUout_F3_2_2  , Final_124_F3_2_2  );
OneRegister RAM_OUT_124_F4_1_1   ( clk , write2_124  , RELUout_F4_1_1  , Final_124_F4_1_1  );
OneRegister RAM_OUT_124_F4_1_2   ( clk , write2_124  , RELUout_F4_1_2  , Final_124_F4_1_2  );
OneRegister RAM_OUT_124_F4_2_1   ( clk , write2_124  , RELUout_F4_2_1  , Final_124_F4_2_1  );
OneRegister RAM_OUT_124_F4_2_2   ( clk , write2_124  , RELUout_F4_2_2  , Final_124_F4_2_2  );
OneRegister RAM_OUT_125_F1_1_1   ( clk , write2_125  , RELUout_F1_1_1  , Final_125_F1_1_1  );
OneRegister RAM_OUT_125_F1_1_2   ( clk , write2_125  , RELUout_F1_1_2  , Final_125_F1_1_2  );
OneRegister RAM_OUT_125_F1_2_1   ( clk , write2_125  , RELUout_F1_2_1  , Final_125_F1_2_1  );
OneRegister RAM_OUT_125_F1_2_2   ( clk , write2_125  , RELUout_F1_2_2  , Final_125_F1_2_2  );
OneRegister RAM_OUT_125_F2_1_1   ( clk , write2_125  , RELUout_F2_1_1  , Final_125_F2_1_1  );
OneRegister RAM_OUT_125_F2_1_2   ( clk , write2_125  , RELUout_F2_1_2  , Final_125_F2_1_2  );
OneRegister RAM_OUT_125_F2_2_1   ( clk , write2_125  , RELUout_F2_2_1  , Final_125_F2_2_1  );
OneRegister RAM_OUT_125_F2_2_2   ( clk , write2_125  , RELUout_F2_2_2  , Final_125_F2_2_2  );
OneRegister RAM_OUT_125_F3_1_1   ( clk , write2_125  , RELUout_F3_1_1  , Final_125_F3_1_1  );
OneRegister RAM_OUT_125_F3_1_2   ( clk , write2_125  , RELUout_F3_1_2  , Final_125_F3_1_2  );
OneRegister RAM_OUT_125_F3_2_1   ( clk , write2_125  , RELUout_F3_2_1  , Final_125_F3_2_1  );
OneRegister RAM_OUT_125_F3_2_2   ( clk , write2_125  , RELUout_F3_2_2  , Final_125_F3_2_2  );
OneRegister RAM_OUT_125_F4_1_1   ( clk , write2_125  , RELUout_F4_1_1  , Final_125_F4_1_1  );
OneRegister RAM_OUT_125_F4_1_2   ( clk , write2_125  , RELUout_F4_1_2  , Final_125_F4_1_2  );
OneRegister RAM_OUT_125_F4_2_1   ( clk , write2_125  , RELUout_F4_2_1  , Final_125_F4_2_1  );
OneRegister RAM_OUT_125_F4_2_2   ( clk , write2_125  , RELUout_F4_2_2  , Final_125_F4_2_2  );
OneRegister RAM_OUT_126_F1_1_1   ( clk , write2_126  , RELUout_F1_1_1  , Final_126_F1_1_1  );
OneRegister RAM_OUT_126_F1_1_2   ( clk , write2_126  , RELUout_F1_1_2  , Final_126_F1_1_2  );
OneRegister RAM_OUT_126_F1_2_1   ( clk , write2_126  , RELUout_F1_2_1  , Final_126_F1_2_1  );
OneRegister RAM_OUT_126_F1_2_2   ( clk , write2_126  , RELUout_F1_2_2  , Final_126_F1_2_2  );
OneRegister RAM_OUT_126_F2_1_1   ( clk , write2_126  , RELUout_F2_1_1  , Final_126_F2_1_1  );
OneRegister RAM_OUT_126_F2_1_2   ( clk , write2_126  , RELUout_F2_1_2  , Final_126_F2_1_2  );
OneRegister RAM_OUT_126_F2_2_1   ( clk , write2_126  , RELUout_F2_2_1  , Final_126_F2_2_1  );
OneRegister RAM_OUT_126_F2_2_2   ( clk , write2_126  , RELUout_F2_2_2  , Final_126_F2_2_2  );
OneRegister RAM_OUT_126_F3_1_1   ( clk , write2_126  , RELUout_F3_1_1  , Final_126_F3_1_1  );
OneRegister RAM_OUT_126_F3_1_2   ( clk , write2_126  , RELUout_F3_1_2  , Final_126_F3_1_2  );
OneRegister RAM_OUT_126_F3_2_1   ( clk , write2_126  , RELUout_F3_2_1  , Final_126_F3_2_1  );
OneRegister RAM_OUT_126_F3_2_2   ( clk , write2_126  , RELUout_F3_2_2  , Final_126_F3_2_2  );
OneRegister RAM_OUT_126_F4_1_1   ( clk , write2_126  , RELUout_F4_1_1  , Final_126_F4_1_1  );
OneRegister RAM_OUT_126_F4_1_2   ( clk , write2_126  , RELUout_F4_1_2  , Final_126_F4_1_2  );
OneRegister RAM_OUT_126_F4_2_1   ( clk , write2_126  , RELUout_F4_2_1  , Final_126_F4_2_1  );
OneRegister RAM_OUT_126_F4_2_2   ( clk , write2_126  , RELUout_F4_2_2  , Final_126_F4_2_2  );
OneRegister RAM_OUT_127_F1_1_1   ( clk , write2_127  , RELUout_F1_1_1  , Final_127_F1_1_1  );
OneRegister RAM_OUT_127_F1_1_2   ( clk , write2_127  , RELUout_F1_1_2  , Final_127_F1_1_2  );
OneRegister RAM_OUT_127_F1_2_1   ( clk , write2_127  , RELUout_F1_2_1  , Final_127_F1_2_1  );
OneRegister RAM_OUT_127_F1_2_2   ( clk , write2_127  , RELUout_F1_2_2  , Final_127_F1_2_2  );
OneRegister RAM_OUT_127_F2_1_1   ( clk , write2_127  , RELUout_F2_1_1  , Final_127_F2_1_1  );
OneRegister RAM_OUT_127_F2_1_2   ( clk , write2_127  , RELUout_F2_1_2  , Final_127_F2_1_2  );
OneRegister RAM_OUT_127_F2_2_1   ( clk , write2_127  , RELUout_F2_2_1  , Final_127_F2_2_1  );
OneRegister RAM_OUT_127_F2_2_2   ( clk , write2_127  , RELUout_F2_2_2  , Final_127_F2_2_2  );
OneRegister RAM_OUT_127_F3_1_1   ( clk , write2_127  , RELUout_F3_1_1  , Final_127_F3_1_1  );
OneRegister RAM_OUT_127_F3_1_2   ( clk , write2_127  , RELUout_F3_1_2  , Final_127_F3_1_2  );
OneRegister RAM_OUT_127_F3_2_1   ( clk , write2_127  , RELUout_F3_2_1  , Final_127_F3_2_1  );
OneRegister RAM_OUT_127_F3_2_2   ( clk , write2_127  , RELUout_F3_2_2  , Final_127_F3_2_2  );
OneRegister RAM_OUT_127_F4_1_1   ( clk , write2_127  , RELUout_F4_1_1  , Final_127_F4_1_1  );
OneRegister RAM_OUT_127_F4_1_2   ( clk , write2_127  , RELUout_F4_1_2  , Final_127_F4_1_2  );
OneRegister RAM_OUT_127_F4_2_1   ( clk , write2_127  , RELUout_F4_2_1  , Final_127_F4_2_1  );
OneRegister RAM_OUT_127_F4_2_2   ( clk , write2_127  , RELUout_F4_2_2  , Final_127_F4_2_2  );
OneRegister RAM_OUT_128_F1_1_1   ( clk , write2_128  , RELUout_F1_1_1  , Final_128_F1_1_1  );
OneRegister RAM_OUT_128_F1_1_2   ( clk , write2_128  , RELUout_F1_1_2  , Final_128_F1_1_2  );
OneRegister RAM_OUT_128_F1_2_1   ( clk , write2_128  , RELUout_F1_2_1  , Final_128_F1_2_1  );
OneRegister RAM_OUT_128_F1_2_2   ( clk , write2_128  , RELUout_F1_2_2  , Final_128_F1_2_2  );
OneRegister RAM_OUT_128_F2_1_1   ( clk , write2_128  , RELUout_F2_1_1  , Final_128_F2_1_1  );
OneRegister RAM_OUT_128_F2_1_2   ( clk , write2_128  , RELUout_F2_1_2  , Final_128_F2_1_2  );
OneRegister RAM_OUT_128_F2_2_1   ( clk , write2_128  , RELUout_F2_2_1  , Final_128_F2_2_1  );
OneRegister RAM_OUT_128_F2_2_2   ( clk , write2_128  , RELUout_F2_2_2  , Final_128_F2_2_2  );
OneRegister RAM_OUT_128_F3_1_1   ( clk , write2_128  , RELUout_F3_1_1  , Final_128_F3_1_1  );
OneRegister RAM_OUT_128_F3_1_2   ( clk , write2_128  , RELUout_F3_1_2  , Final_128_F3_1_2  );
OneRegister RAM_OUT_128_F3_2_1   ( clk , write2_128  , RELUout_F3_2_1  , Final_128_F3_2_1  );
OneRegister RAM_OUT_128_F3_2_2   ( clk , write2_128  , RELUout_F3_2_2  , Final_128_F3_2_2  );
OneRegister RAM_OUT_128_F4_1_1   ( clk , write2_128  , RELUout_F4_1_1  , Final_128_F4_1_1  );
OneRegister RAM_OUT_128_F4_1_2   ( clk , write2_128  , RELUout_F4_1_2  , Final_128_F4_1_2  );
OneRegister RAM_OUT_128_F4_2_1   ( clk , write2_128  , RELUout_F4_2_1  , Final_128_F4_2_1  );
OneRegister RAM_OUT_128_F4_2_2   ( clk , write2_128  , RELUout_F4_2_2  , Final_128_F4_2_2  );
OneRegister RAM_OUT_129_F1_1_1   ( clk , write2_129  , RELUout_F1_1_1  , Final_129_F1_1_1  );
OneRegister RAM_OUT_129_F1_1_2   ( clk , write2_129  , RELUout_F1_1_2  , Final_129_F1_1_2  );
OneRegister RAM_OUT_129_F1_2_1   ( clk , write2_129  , RELUout_F1_2_1  , Final_129_F1_2_1  );
OneRegister RAM_OUT_129_F1_2_2   ( clk , write2_129  , RELUout_F1_2_2  , Final_129_F1_2_2  );
OneRegister RAM_OUT_129_F2_1_1   ( clk , write2_129  , RELUout_F2_1_1  , Final_129_F2_1_1  );
OneRegister RAM_OUT_129_F2_1_2   ( clk , write2_129  , RELUout_F2_1_2  , Final_129_F2_1_2  );
OneRegister RAM_OUT_129_F2_2_1   ( clk , write2_129  , RELUout_F2_2_1  , Final_129_F2_2_1  );
OneRegister RAM_OUT_129_F2_2_2   ( clk , write2_129  , RELUout_F2_2_2  , Final_129_F2_2_2  );
OneRegister RAM_OUT_129_F3_1_1   ( clk , write2_129  , RELUout_F3_1_1  , Final_129_F3_1_1  );
OneRegister RAM_OUT_129_F3_1_2   ( clk , write2_129  , RELUout_F3_1_2  , Final_129_F3_1_2  );
OneRegister RAM_OUT_129_F3_2_1   ( clk , write2_129  , RELUout_F3_2_1  , Final_129_F3_2_1  );
OneRegister RAM_OUT_129_F3_2_2   ( clk , write2_129  , RELUout_F3_2_2  , Final_129_F3_2_2  );
OneRegister RAM_OUT_129_F4_1_1   ( clk , write2_129  , RELUout_F4_1_1  , Final_129_F4_1_1  );
OneRegister RAM_OUT_129_F4_1_2   ( clk , write2_129  , RELUout_F4_1_2  , Final_129_F4_1_2  );
OneRegister RAM_OUT_129_F4_2_1   ( clk , write2_129  , RELUout_F4_2_1  , Final_129_F4_2_1  );
OneRegister RAM_OUT_129_F4_2_2   ( clk , write2_129  , RELUout_F4_2_2  , Final_129_F4_2_2  );
OneRegister RAM_OUT_130_F1_1_1   ( clk , write2_130  , RELUout_F1_1_1  , Final_130_F1_1_1  );
OneRegister RAM_OUT_130_F1_1_2   ( clk , write2_130  , RELUout_F1_1_2  , Final_130_F1_1_2  );
OneRegister RAM_OUT_130_F1_2_1   ( clk , write2_130  , RELUout_F1_2_1  , Final_130_F1_2_1  );
OneRegister RAM_OUT_130_F1_2_2   ( clk , write2_130  , RELUout_F1_2_2  , Final_130_F1_2_2  );
OneRegister RAM_OUT_130_F2_1_1   ( clk , write2_130  , RELUout_F2_1_1  , Final_130_F2_1_1  );
OneRegister RAM_OUT_130_F2_1_2   ( clk , write2_130  , RELUout_F2_1_2  , Final_130_F2_1_2  );
OneRegister RAM_OUT_130_F2_2_1   ( clk , write2_130  , RELUout_F2_2_1  , Final_130_F2_2_1  );
OneRegister RAM_OUT_130_F2_2_2   ( clk , write2_130  , RELUout_F2_2_2  , Final_130_F2_2_2  );
OneRegister RAM_OUT_130_F3_1_1   ( clk , write2_130  , RELUout_F3_1_1  , Final_130_F3_1_1  );
OneRegister RAM_OUT_130_F3_1_2   ( clk , write2_130  , RELUout_F3_1_2  , Final_130_F3_1_2  );
OneRegister RAM_OUT_130_F3_2_1   ( clk , write2_130  , RELUout_F3_2_1  , Final_130_F3_2_1  );
OneRegister RAM_OUT_130_F3_2_2   ( clk , write2_130  , RELUout_F3_2_2  , Final_130_F3_2_2  );
OneRegister RAM_OUT_130_F4_1_1   ( clk , write2_130  , RELUout_F4_1_1  , Final_130_F4_1_1  );
OneRegister RAM_OUT_130_F4_1_2   ( clk , write2_130  , RELUout_F4_1_2  , Final_130_F4_1_2  );
OneRegister RAM_OUT_130_F4_2_1   ( clk , write2_130  , RELUout_F4_2_1  , Final_130_F4_2_1  );
OneRegister RAM_OUT_130_F4_2_2   ( clk , write2_130  , RELUout_F4_2_2  , Final_130_F4_2_2  );
OneRegister RAM_OUT_131_F1_1_1   ( clk , write2_131  , RELUout_F1_1_1  , Final_131_F1_1_1  );
OneRegister RAM_OUT_131_F1_1_2   ( clk , write2_131  , RELUout_F1_1_2  , Final_131_F1_1_2  );
OneRegister RAM_OUT_131_F1_2_1   ( clk , write2_131  , RELUout_F1_2_1  , Final_131_F1_2_1  );
OneRegister RAM_OUT_131_F1_2_2   ( clk , write2_131  , RELUout_F1_2_2  , Final_131_F1_2_2  );
OneRegister RAM_OUT_131_F2_1_1   ( clk , write2_131  , RELUout_F2_1_1  , Final_131_F2_1_1  );
OneRegister RAM_OUT_131_F2_1_2   ( clk , write2_131  , RELUout_F2_1_2  , Final_131_F2_1_2  );
OneRegister RAM_OUT_131_F2_2_1   ( clk , write2_131  , RELUout_F2_2_1  , Final_131_F2_2_1  );
OneRegister RAM_OUT_131_F2_2_2   ( clk , write2_131  , RELUout_F2_2_2  , Final_131_F2_2_2  );
OneRegister RAM_OUT_131_F3_1_1   ( clk , write2_131  , RELUout_F3_1_1  , Final_131_F3_1_1  );
OneRegister RAM_OUT_131_F3_1_2   ( clk , write2_131  , RELUout_F3_1_2  , Final_131_F3_1_2  );
OneRegister RAM_OUT_131_F3_2_1   ( clk , write2_131  , RELUout_F3_2_1  , Final_131_F3_2_1  );
OneRegister RAM_OUT_131_F3_2_2   ( clk , write2_131  , RELUout_F3_2_2  , Final_131_F3_2_2  );
OneRegister RAM_OUT_131_F4_1_1   ( clk , write2_131  , RELUout_F4_1_1  , Final_131_F4_1_1  );
OneRegister RAM_OUT_131_F4_1_2   ( clk , write2_131  , RELUout_F4_1_2  , Final_131_F4_1_2  );
OneRegister RAM_OUT_131_F4_2_1   ( clk , write2_131  , RELUout_F4_2_1  , Final_131_F4_2_1  );
OneRegister RAM_OUT_131_F4_2_2   ( clk , write2_131  , RELUout_F4_2_2  , Final_131_F4_2_2  );
OneRegister RAM_OUT_132_F1_1_1   ( clk , write2_132  , RELUout_F1_1_1  , Final_132_F1_1_1  );
OneRegister RAM_OUT_132_F1_1_2   ( clk , write2_132  , RELUout_F1_1_2  , Final_132_F1_1_2  );
OneRegister RAM_OUT_132_F1_2_1   ( clk , write2_132  , RELUout_F1_2_1  , Final_132_F1_2_1  );
OneRegister RAM_OUT_132_F1_2_2   ( clk , write2_132  , RELUout_F1_2_2  , Final_132_F1_2_2  );
OneRegister RAM_OUT_132_F2_1_1   ( clk , write2_132  , RELUout_F2_1_1  , Final_132_F2_1_1  );
OneRegister RAM_OUT_132_F2_1_2   ( clk , write2_132  , RELUout_F2_1_2  , Final_132_F2_1_2  );
OneRegister RAM_OUT_132_F2_2_1   ( clk , write2_132  , RELUout_F2_2_1  , Final_132_F2_2_1  );
OneRegister RAM_OUT_132_F2_2_2   ( clk , write2_132  , RELUout_F2_2_2  , Final_132_F2_2_2  );
OneRegister RAM_OUT_132_F3_1_1   ( clk , write2_132  , RELUout_F3_1_1  , Final_132_F3_1_1  );
OneRegister RAM_OUT_132_F3_1_2   ( clk , write2_132  , RELUout_F3_1_2  , Final_132_F3_1_2  );
OneRegister RAM_OUT_132_F3_2_1   ( clk , write2_132  , RELUout_F3_2_1  , Final_132_F3_2_1  );
OneRegister RAM_OUT_132_F3_2_2   ( clk , write2_132  , RELUout_F3_2_2  , Final_132_F3_2_2  );
OneRegister RAM_OUT_132_F4_1_1   ( clk , write2_132  , RELUout_F4_1_1  , Final_132_F4_1_1  );
OneRegister RAM_OUT_132_F4_1_2   ( clk , write2_132  , RELUout_F4_1_2  , Final_132_F4_1_2  );
OneRegister RAM_OUT_132_F4_2_1   ( clk , write2_132  , RELUout_F4_2_1  , Final_132_F4_2_1  );
OneRegister RAM_OUT_132_F4_2_2   ( clk , write2_132  , RELUout_F4_2_2  , Final_132_F4_2_2  );
OneRegister RAM_OUT_133_F1_1_1   ( clk , write2_133  , RELUout_F1_1_1  , Final_133_F1_1_1  );
OneRegister RAM_OUT_133_F1_1_2   ( clk , write2_133  , RELUout_F1_1_2  , Final_133_F1_1_2  );
OneRegister RAM_OUT_133_F1_2_1   ( clk , write2_133  , RELUout_F1_2_1  , Final_133_F1_2_1  );
OneRegister RAM_OUT_133_F1_2_2   ( clk , write2_133  , RELUout_F1_2_2  , Final_133_F1_2_2  );
OneRegister RAM_OUT_133_F2_1_1   ( clk , write2_133  , RELUout_F2_1_1  , Final_133_F2_1_1  );
OneRegister RAM_OUT_133_F2_1_2   ( clk , write2_133  , RELUout_F2_1_2  , Final_133_F2_1_2  );
OneRegister RAM_OUT_133_F2_2_1   ( clk , write2_133  , RELUout_F2_2_1  , Final_133_F2_2_1  );
OneRegister RAM_OUT_133_F2_2_2   ( clk , write2_133  , RELUout_F2_2_2  , Final_133_F2_2_2  );
OneRegister RAM_OUT_133_F3_1_1   ( clk , write2_133  , RELUout_F3_1_1  , Final_133_F3_1_1  );
OneRegister RAM_OUT_133_F3_1_2   ( clk , write2_133  , RELUout_F3_1_2  , Final_133_F3_1_2  );
OneRegister RAM_OUT_133_F3_2_1   ( clk , write2_133  , RELUout_F3_2_1  , Final_133_F3_2_1  );
OneRegister RAM_OUT_133_F3_2_2   ( clk , write2_133  , RELUout_F3_2_2  , Final_133_F3_2_2  );
OneRegister RAM_OUT_133_F4_1_1   ( clk , write2_133  , RELUout_F4_1_1  , Final_133_F4_1_1  );
OneRegister RAM_OUT_133_F4_1_2   ( clk , write2_133  , RELUout_F4_1_2  , Final_133_F4_1_2  );
OneRegister RAM_OUT_133_F4_2_1   ( clk , write2_133  , RELUout_F4_2_1  , Final_133_F4_2_1  );
OneRegister RAM_OUT_133_F4_2_2   ( clk , write2_133  , RELUout_F4_2_2  , Final_133_F4_2_2  );
OneRegister RAM_OUT_134_F1_1_1   ( clk , write2_134  , RELUout_F1_1_1  , Final_134_F1_1_1  );
OneRegister RAM_OUT_134_F1_1_2   ( clk , write2_134  , RELUout_F1_1_2  , Final_134_F1_1_2  );
OneRegister RAM_OUT_134_F1_2_1   ( clk , write2_134  , RELUout_F1_2_1  , Final_134_F1_2_1  );
OneRegister RAM_OUT_134_F1_2_2   ( clk , write2_134  , RELUout_F1_2_2  , Final_134_F1_2_2  );
OneRegister RAM_OUT_134_F2_1_1   ( clk , write2_134  , RELUout_F2_1_1  , Final_134_F2_1_1  );
OneRegister RAM_OUT_134_F2_1_2   ( clk , write2_134  , RELUout_F2_1_2  , Final_134_F2_1_2  );
OneRegister RAM_OUT_134_F2_2_1   ( clk , write2_134  , RELUout_F2_2_1  , Final_134_F2_2_1  );
OneRegister RAM_OUT_134_F2_2_2   ( clk , write2_134  , RELUout_F2_2_2  , Final_134_F2_2_2  );
OneRegister RAM_OUT_134_F3_1_1   ( clk , write2_134  , RELUout_F3_1_1  , Final_134_F3_1_1  );
OneRegister RAM_OUT_134_F3_1_2   ( clk , write2_134  , RELUout_F3_1_2  , Final_134_F3_1_2  );
OneRegister RAM_OUT_134_F3_2_1   ( clk , write2_134  , RELUout_F3_2_1  , Final_134_F3_2_1  );
OneRegister RAM_OUT_134_F3_2_2   ( clk , write2_134  , RELUout_F3_2_2  , Final_134_F3_2_2  );
OneRegister RAM_OUT_134_F4_1_1   ( clk , write2_134  , RELUout_F4_1_1  , Final_134_F4_1_1  );
OneRegister RAM_OUT_134_F4_1_2   ( clk , write2_134  , RELUout_F4_1_2  , Final_134_F4_1_2  );
OneRegister RAM_OUT_134_F4_2_1   ( clk , write2_134  , RELUout_F4_2_1  , Final_134_F4_2_1  );
OneRegister RAM_OUT_134_F4_2_2   ( clk , write2_134  , RELUout_F4_2_2  , Final_134_F4_2_2  );
OneRegister RAM_OUT_135_F1_1_1   ( clk , write2_135  , RELUout_F1_1_1  , Final_135_F1_1_1  );
OneRegister RAM_OUT_135_F1_1_2   ( clk , write2_135  , RELUout_F1_1_2  , Final_135_F1_1_2  );
OneRegister RAM_OUT_135_F1_2_1   ( clk , write2_135  , RELUout_F1_2_1  , Final_135_F1_2_1  );
OneRegister RAM_OUT_135_F1_2_2   ( clk , write2_135  , RELUout_F1_2_2  , Final_135_F1_2_2  );
OneRegister RAM_OUT_135_F2_1_1   ( clk , write2_135  , RELUout_F2_1_1  , Final_135_F2_1_1  );
OneRegister RAM_OUT_135_F2_1_2   ( clk , write2_135  , RELUout_F2_1_2  , Final_135_F2_1_2  );
OneRegister RAM_OUT_135_F2_2_1   ( clk , write2_135  , RELUout_F2_2_1  , Final_135_F2_2_1  );
OneRegister RAM_OUT_135_F2_2_2   ( clk , write2_135  , RELUout_F2_2_2  , Final_135_F2_2_2  );
OneRegister RAM_OUT_135_F3_1_1   ( clk , write2_135  , RELUout_F3_1_1  , Final_135_F3_1_1  );
OneRegister RAM_OUT_135_F3_1_2   ( clk , write2_135  , RELUout_F3_1_2  , Final_135_F3_1_2  );
OneRegister RAM_OUT_135_F3_2_1   ( clk , write2_135  , RELUout_F3_2_1  , Final_135_F3_2_1  );
OneRegister RAM_OUT_135_F3_2_2   ( clk , write2_135  , RELUout_F3_2_2  , Final_135_F3_2_2  );
OneRegister RAM_OUT_135_F4_1_1   ( clk , write2_135  , RELUout_F4_1_1  , Final_135_F4_1_1  );
OneRegister RAM_OUT_135_F4_1_2   ( clk , write2_135  , RELUout_F4_1_2  , Final_135_F4_1_2  );
OneRegister RAM_OUT_135_F4_2_1   ( clk , write2_135  , RELUout_F4_2_1  , Final_135_F4_2_1  );
OneRegister RAM_OUT_135_F4_2_2   ( clk , write2_135  , RELUout_F4_2_2  , Final_135_F4_2_2  );
OneRegister RAM_OUT_136_F1_1_1   ( clk , write2_136  , RELUout_F1_1_1  , Final_136_F1_1_1  );
OneRegister RAM_OUT_136_F1_1_2   ( clk , write2_136  , RELUout_F1_1_2  , Final_136_F1_1_2  );
OneRegister RAM_OUT_136_F1_2_1   ( clk , write2_136  , RELUout_F1_2_1  , Final_136_F1_2_1  );
OneRegister RAM_OUT_136_F1_2_2   ( clk , write2_136  , RELUout_F1_2_2  , Final_136_F1_2_2  );
OneRegister RAM_OUT_136_F2_1_1   ( clk , write2_136  , RELUout_F2_1_1  , Final_136_F2_1_1  );
OneRegister RAM_OUT_136_F2_1_2   ( clk , write2_136  , RELUout_F2_1_2  , Final_136_F2_1_2  );
OneRegister RAM_OUT_136_F2_2_1   ( clk , write2_136  , RELUout_F2_2_1  , Final_136_F2_2_1  );
OneRegister RAM_OUT_136_F2_2_2   ( clk , write2_136  , RELUout_F2_2_2  , Final_136_F2_2_2  );
OneRegister RAM_OUT_136_F3_1_1   ( clk , write2_136  , RELUout_F3_1_1  , Final_136_F3_1_1  );
OneRegister RAM_OUT_136_F3_1_2   ( clk , write2_136  , RELUout_F3_1_2  , Final_136_F3_1_2  );
OneRegister RAM_OUT_136_F3_2_1   ( clk , write2_136  , RELUout_F3_2_1  , Final_136_F3_2_1  );
OneRegister RAM_OUT_136_F3_2_2   ( clk , write2_136  , RELUout_F3_2_2  , Final_136_F3_2_2  );
OneRegister RAM_OUT_136_F4_1_1   ( clk , write2_136  , RELUout_F4_1_1  , Final_136_F4_1_1  );
OneRegister RAM_OUT_136_F4_1_2   ( clk , write2_136  , RELUout_F4_1_2  , Final_136_F4_1_2  );
OneRegister RAM_OUT_136_F4_2_1   ( clk , write2_136  , RELUout_F4_2_1  , Final_136_F4_2_1  );
OneRegister RAM_OUT_136_F4_2_2   ( clk , write2_136  , RELUout_F4_2_2  , Final_136_F4_2_2  );
OneRegister RAM_OUT_137_F1_1_1   ( clk , write2_137  , RELUout_F1_1_1  , Final_137_F1_1_1  );
OneRegister RAM_OUT_137_F1_1_2   ( clk , write2_137  , RELUout_F1_1_2  , Final_137_F1_1_2  );
OneRegister RAM_OUT_137_F1_2_1   ( clk , write2_137  , RELUout_F1_2_1  , Final_137_F1_2_1  );
OneRegister RAM_OUT_137_F1_2_2   ( clk , write2_137  , RELUout_F1_2_2  , Final_137_F1_2_2  );
OneRegister RAM_OUT_137_F2_1_1   ( clk , write2_137  , RELUout_F2_1_1  , Final_137_F2_1_1  );
OneRegister RAM_OUT_137_F2_1_2   ( clk , write2_137  , RELUout_F2_1_2  , Final_137_F2_1_2  );
OneRegister RAM_OUT_137_F2_2_1   ( clk , write2_137  , RELUout_F2_2_1  , Final_137_F2_2_1  );
OneRegister RAM_OUT_137_F2_2_2   ( clk , write2_137  , RELUout_F2_2_2  , Final_137_F2_2_2  );
OneRegister RAM_OUT_137_F3_1_1   ( clk , write2_137  , RELUout_F3_1_1  , Final_137_F3_1_1  );
OneRegister RAM_OUT_137_F3_1_2   ( clk , write2_137  , RELUout_F3_1_2  , Final_137_F3_1_2  );
OneRegister RAM_OUT_137_F3_2_1   ( clk , write2_137  , RELUout_F3_2_1  , Final_137_F3_2_1  );
OneRegister RAM_OUT_137_F3_2_2   ( clk , write2_137  , RELUout_F3_2_2  , Final_137_F3_2_2  );
OneRegister RAM_OUT_137_F4_1_1   ( clk , write2_137  , RELUout_F4_1_1  , Final_137_F4_1_1  );
OneRegister RAM_OUT_137_F4_1_2   ( clk , write2_137  , RELUout_F4_1_2  , Final_137_F4_1_2  );
OneRegister RAM_OUT_137_F4_2_1   ( clk , write2_137  , RELUout_F4_2_1  , Final_137_F4_2_1  );
OneRegister RAM_OUT_137_F4_2_2   ( clk , write2_137  , RELUout_F4_2_2  , Final_137_F4_2_2  );
OneRegister RAM_OUT_138_F1_1_1   ( clk , write2_138  , RELUout_F1_1_1  , Final_138_F1_1_1  );
OneRegister RAM_OUT_138_F1_1_2   ( clk , write2_138  , RELUout_F1_1_2  , Final_138_F1_1_2  );
OneRegister RAM_OUT_138_F1_2_1   ( clk , write2_138  , RELUout_F1_2_1  , Final_138_F1_2_1  );
OneRegister RAM_OUT_138_F1_2_2   ( clk , write2_138  , RELUout_F1_2_2  , Final_138_F1_2_2  );
OneRegister RAM_OUT_138_F2_1_1   ( clk , write2_138  , RELUout_F2_1_1  , Final_138_F2_1_1  );
OneRegister RAM_OUT_138_F2_1_2   ( clk , write2_138  , RELUout_F2_1_2  , Final_138_F2_1_2  );
OneRegister RAM_OUT_138_F2_2_1   ( clk , write2_138  , RELUout_F2_2_1  , Final_138_F2_2_1  );
OneRegister RAM_OUT_138_F2_2_2   ( clk , write2_138  , RELUout_F2_2_2  , Final_138_F2_2_2  );
OneRegister RAM_OUT_138_F3_1_1   ( clk , write2_138  , RELUout_F3_1_1  , Final_138_F3_1_1  );
OneRegister RAM_OUT_138_F3_1_2   ( clk , write2_138  , RELUout_F3_1_2  , Final_138_F3_1_2  );
OneRegister RAM_OUT_138_F3_2_1   ( clk , write2_138  , RELUout_F3_2_1  , Final_138_F3_2_1  );
OneRegister RAM_OUT_138_F3_2_2   ( clk , write2_138  , RELUout_F3_2_2  , Final_138_F3_2_2  );
OneRegister RAM_OUT_138_F4_1_1   ( clk , write2_138  , RELUout_F4_1_1  , Final_138_F4_1_1  );
OneRegister RAM_OUT_138_F4_1_2   ( clk , write2_138  , RELUout_F4_1_2  , Final_138_F4_1_2  );
OneRegister RAM_OUT_138_F4_2_1   ( clk , write2_138  , RELUout_F4_2_1  , Final_138_F4_2_1  );
OneRegister RAM_OUT_138_F4_2_2   ( clk , write2_138  , RELUout_F4_2_2  , Final_138_F4_2_2  );
OneRegister RAM_OUT_139_F1_1_1   ( clk , write2_139  , RELUout_F1_1_1  , Final_139_F1_1_1  );
OneRegister RAM_OUT_139_F1_1_2   ( clk , write2_139  , RELUout_F1_1_2  , Final_139_F1_1_2  );
OneRegister RAM_OUT_139_F1_2_1   ( clk , write2_139  , RELUout_F1_2_1  , Final_139_F1_2_1  );
OneRegister RAM_OUT_139_F1_2_2   ( clk , write2_139  , RELUout_F1_2_2  , Final_139_F1_2_2  );
OneRegister RAM_OUT_139_F2_1_1   ( clk , write2_139  , RELUout_F2_1_1  , Final_139_F2_1_1  );
OneRegister RAM_OUT_139_F2_1_2   ( clk , write2_139  , RELUout_F2_1_2  , Final_139_F2_1_2  );
OneRegister RAM_OUT_139_F2_2_1   ( clk , write2_139  , RELUout_F2_2_1  , Final_139_F2_2_1  );
OneRegister RAM_OUT_139_F2_2_2   ( clk , write2_139  , RELUout_F2_2_2  , Final_139_F2_2_2  );
OneRegister RAM_OUT_139_F3_1_1   ( clk , write2_139  , RELUout_F3_1_1  , Final_139_F3_1_1  );
OneRegister RAM_OUT_139_F3_1_2   ( clk , write2_139  , RELUout_F3_1_2  , Final_139_F3_1_2  );
OneRegister RAM_OUT_139_F3_2_1   ( clk , write2_139  , RELUout_F3_2_1  , Final_139_F3_2_1  );
OneRegister RAM_OUT_139_F3_2_2   ( clk , write2_139  , RELUout_F3_2_2  , Final_139_F3_2_2  );
OneRegister RAM_OUT_139_F4_1_1   ( clk , write2_139  , RELUout_F4_1_1  , Final_139_F4_1_1  );
OneRegister RAM_OUT_139_F4_1_2   ( clk , write2_139  , RELUout_F4_1_2  , Final_139_F4_1_2  );
OneRegister RAM_OUT_139_F4_2_1   ( clk , write2_139  , RELUout_F4_2_1  , Final_139_F4_2_1  );
OneRegister RAM_OUT_139_F4_2_2   ( clk , write2_139  , RELUout_F4_2_2  , Final_139_F4_2_2  );
OneRegister RAM_OUT_140_F1_1_1   ( clk , write2_140  , RELUout_F1_1_1  , Final_140_F1_1_1  );
OneRegister RAM_OUT_140_F1_1_2   ( clk , write2_140  , RELUout_F1_1_2  , Final_140_F1_1_2  );
OneRegister RAM_OUT_140_F1_2_1   ( clk , write2_140  , RELUout_F1_2_1  , Final_140_F1_2_1  );
OneRegister RAM_OUT_140_F1_2_2   ( clk , write2_140  , RELUout_F1_2_2  , Final_140_F1_2_2  );
OneRegister RAM_OUT_140_F2_1_1   ( clk , write2_140  , RELUout_F2_1_1  , Final_140_F2_1_1  );
OneRegister RAM_OUT_140_F2_1_2   ( clk , write2_140  , RELUout_F2_1_2  , Final_140_F2_1_2  );
OneRegister RAM_OUT_140_F2_2_1   ( clk , write2_140  , RELUout_F2_2_1  , Final_140_F2_2_1  );
OneRegister RAM_OUT_140_F2_2_2   ( clk , write2_140  , RELUout_F2_2_2  , Final_140_F2_2_2  );
OneRegister RAM_OUT_140_F3_1_1   ( clk , write2_140  , RELUout_F3_1_1  , Final_140_F3_1_1  );
OneRegister RAM_OUT_140_F3_1_2   ( clk , write2_140  , RELUout_F3_1_2  , Final_140_F3_1_2  );
OneRegister RAM_OUT_140_F3_2_1   ( clk , write2_140  , RELUout_F3_2_1  , Final_140_F3_2_1  );
OneRegister RAM_OUT_140_F3_2_2   ( clk , write2_140  , RELUout_F3_2_2  , Final_140_F3_2_2  );
OneRegister RAM_OUT_140_F4_1_1   ( clk , write2_140  , RELUout_F4_1_1  , Final_140_F4_1_1  );
OneRegister RAM_OUT_140_F4_1_2   ( clk , write2_140  , RELUout_F4_1_2  , Final_140_F4_1_2  );
OneRegister RAM_OUT_140_F4_2_1   ( clk , write2_140  , RELUout_F4_2_1  , Final_140_F4_2_1  );
OneRegister RAM_OUT_140_F4_2_2   ( clk , write2_140  , RELUout_F4_2_2  , Final_140_F4_2_2  );
OneRegister RAM_OUT_141_F1_1_1   ( clk , write2_141  , RELUout_F1_1_1  , Final_141_F1_1_1  );
OneRegister RAM_OUT_141_F1_1_2   ( clk , write2_141  , RELUout_F1_1_2  , Final_141_F1_1_2  );
OneRegister RAM_OUT_141_F1_2_1   ( clk , write2_141  , RELUout_F1_2_1  , Final_141_F1_2_1  );
OneRegister RAM_OUT_141_F1_2_2   ( clk , write2_141  , RELUout_F1_2_2  , Final_141_F1_2_2  );
OneRegister RAM_OUT_141_F2_1_1   ( clk , write2_141  , RELUout_F2_1_1  , Final_141_F2_1_1  );
OneRegister RAM_OUT_141_F2_1_2   ( clk , write2_141  , RELUout_F2_1_2  , Final_141_F2_1_2  );
OneRegister RAM_OUT_141_F2_2_1   ( clk , write2_141  , RELUout_F2_2_1  , Final_141_F2_2_1  );
OneRegister RAM_OUT_141_F2_2_2   ( clk , write2_141  , RELUout_F2_2_2  , Final_141_F2_2_2  );
OneRegister RAM_OUT_141_F3_1_1   ( clk , write2_141  , RELUout_F3_1_1  , Final_141_F3_1_1  );
OneRegister RAM_OUT_141_F3_1_2   ( clk , write2_141  , RELUout_F3_1_2  , Final_141_F3_1_2  );
OneRegister RAM_OUT_141_F3_2_1   ( clk , write2_141  , RELUout_F3_2_1  , Final_141_F3_2_1  );
OneRegister RAM_OUT_141_F3_2_2   ( clk , write2_141  , RELUout_F3_2_2  , Final_141_F3_2_2  );
OneRegister RAM_OUT_141_F4_1_1   ( clk , write2_141  , RELUout_F4_1_1  , Final_141_F4_1_1  );
OneRegister RAM_OUT_141_F4_1_2   ( clk , write2_141  , RELUout_F4_1_2  , Final_141_F4_1_2  );
OneRegister RAM_OUT_141_F4_2_1   ( clk , write2_141  , RELUout_F4_2_1  , Final_141_F4_2_1  );
OneRegister RAM_OUT_141_F4_2_2   ( clk , write2_141  , RELUout_F4_2_2  , Final_141_F4_2_2  );
OneRegister RAM_OUT_142_F1_1_1   ( clk , write2_142  , RELUout_F1_1_1  , Final_142_F1_1_1  );
OneRegister RAM_OUT_142_F1_1_2   ( clk , write2_142  , RELUout_F1_1_2  , Final_142_F1_1_2  );
OneRegister RAM_OUT_142_F1_2_1   ( clk , write2_142  , RELUout_F1_2_1  , Final_142_F1_2_1  );
OneRegister RAM_OUT_142_F1_2_2   ( clk , write2_142  , RELUout_F1_2_2  , Final_142_F1_2_2  );
OneRegister RAM_OUT_142_F2_1_1   ( clk , write2_142  , RELUout_F2_1_1  , Final_142_F2_1_1  );
OneRegister RAM_OUT_142_F2_1_2   ( clk , write2_142  , RELUout_F2_1_2  , Final_142_F2_1_2  );
OneRegister RAM_OUT_142_F2_2_1   ( clk , write2_142  , RELUout_F2_2_1  , Final_142_F2_2_1  );
OneRegister RAM_OUT_142_F2_2_2   ( clk , write2_142  , RELUout_F2_2_2  , Final_142_F2_2_2  );
OneRegister RAM_OUT_142_F3_1_1   ( clk , write2_142  , RELUout_F3_1_1  , Final_142_F3_1_1  );
OneRegister RAM_OUT_142_F3_1_2   ( clk , write2_142  , RELUout_F3_1_2  , Final_142_F3_1_2  );
OneRegister RAM_OUT_142_F3_2_1   ( clk , write2_142  , RELUout_F3_2_1  , Final_142_F3_2_1  );
OneRegister RAM_OUT_142_F3_2_2   ( clk , write2_142  , RELUout_F3_2_2  , Final_142_F3_2_2  );
OneRegister RAM_OUT_142_F4_1_1   ( clk , write2_142  , RELUout_F4_1_1  , Final_142_F4_1_1  );
OneRegister RAM_OUT_142_F4_1_2   ( clk , write2_142  , RELUout_F4_1_2  , Final_142_F4_1_2  );
OneRegister RAM_OUT_142_F4_2_1   ( clk , write2_142  , RELUout_F4_2_1  , Final_142_F4_2_1  );
OneRegister RAM_OUT_142_F4_2_2   ( clk , write2_142  , RELUout_F4_2_2  , Final_142_F4_2_2  );
OneRegister RAM_OUT_143_F1_1_1   ( clk , write2_143  , RELUout_F1_1_1  , Final_143_F1_1_1  );
OneRegister RAM_OUT_143_F1_1_2   ( clk , write2_143  , RELUout_F1_1_2  , Final_143_F1_1_2  );
OneRegister RAM_OUT_143_F1_2_1   ( clk , write2_143  , RELUout_F1_2_1  , Final_143_F1_2_1  );
OneRegister RAM_OUT_143_F1_2_2   ( clk , write2_143  , RELUout_F1_2_2  , Final_143_F1_2_2  );
OneRegister RAM_OUT_143_F2_1_1   ( clk , write2_143  , RELUout_F2_1_1  , Final_143_F2_1_1  );
OneRegister RAM_OUT_143_F2_1_2   ( clk , write2_143  , RELUout_F2_1_2  , Final_143_F2_1_2  );
OneRegister RAM_OUT_143_F2_2_1   ( clk , write2_143  , RELUout_F2_2_1  , Final_143_F2_2_1  );
OneRegister RAM_OUT_143_F2_2_2   ( clk , write2_143  , RELUout_F2_2_2  , Final_143_F2_2_2  );
OneRegister RAM_OUT_143_F3_1_1   ( clk , write2_143  , RELUout_F3_1_1  , Final_143_F3_1_1  );
OneRegister RAM_OUT_143_F3_1_2   ( clk , write2_143  , RELUout_F3_1_2  , Final_143_F3_1_2  );
OneRegister RAM_OUT_143_F3_2_1   ( clk , write2_143  , RELUout_F3_2_1  , Final_143_F3_2_1  );
OneRegister RAM_OUT_143_F3_2_2   ( clk , write2_143  , RELUout_F3_2_2  , Final_143_F3_2_2  );
OneRegister RAM_OUT_143_F4_1_1   ( clk , write2_143  , RELUout_F4_1_1  , Final_143_F4_1_1  );
OneRegister RAM_OUT_143_F4_1_2   ( clk , write2_143  , RELUout_F4_1_2  , Final_143_F4_1_2  );
OneRegister RAM_OUT_143_F4_2_1   ( clk , write2_143  , RELUout_F4_2_1  , Final_143_F4_2_1  );
OneRegister RAM_OUT_143_F4_2_2   ( clk , write2_143  , RELUout_F4_2_2  , Final_143_F4_2_2  );
OneRegister RAM_OUT_144_F1_1_1   ( clk , write2_144  , RELUout_F1_1_1  , Final_144_F1_1_1  );
OneRegister RAM_OUT_144_F1_1_2   ( clk , write2_144  , RELUout_F1_1_2  , Final_144_F1_1_2  );
OneRegister RAM_OUT_144_F1_2_1   ( clk , write2_144  , RELUout_F1_2_1  , Final_144_F1_2_1  );
OneRegister RAM_OUT_144_F1_2_2   ( clk , write2_144  , RELUout_F1_2_2  , Final_144_F1_2_2  );
OneRegister RAM_OUT_144_F2_1_1   ( clk , write2_144  , RELUout_F2_1_1  , Final_144_F2_1_1  );
OneRegister RAM_OUT_144_F2_1_2   ( clk , write2_144  , RELUout_F2_1_2  , Final_144_F2_1_2  );
OneRegister RAM_OUT_144_F2_2_1   ( clk , write2_144  , RELUout_F2_2_1  , Final_144_F2_2_1  );
OneRegister RAM_OUT_144_F2_2_2   ( clk , write2_144  , RELUout_F2_2_2  , Final_144_F2_2_2  );
OneRegister RAM_OUT_144_F3_1_1   ( clk , write2_144  , RELUout_F3_1_1  , Final_144_F3_1_1  );
OneRegister RAM_OUT_144_F3_1_2   ( clk , write2_144  , RELUout_F3_1_2  , Final_144_F3_1_2  );
OneRegister RAM_OUT_144_F3_2_1   ( clk , write2_144  , RELUout_F3_2_1  , Final_144_F3_2_1  );
OneRegister RAM_OUT_144_F3_2_2   ( clk , write2_144  , RELUout_F3_2_2  , Final_144_F3_2_2  );
OneRegister RAM_OUT_144_F4_1_1   ( clk , write2_144  , RELUout_F4_1_1  , Final_144_F4_1_1  );
OneRegister RAM_OUT_144_F4_1_2   ( clk , write2_144  , RELUout_F4_1_2  , Final_144_F4_1_2  );
OneRegister RAM_OUT_144_F4_2_1   ( clk , write2_144  , RELUout_F4_2_1  , Final_144_F4_2_1  );
OneRegister RAM_OUT_144_F4_2_2   ( clk , write2_144  , RELUout_F4_2_2  , Final_144_F4_2_2  );

*/

/* endmodule


module MAX1LAYER_bla2_2by2(clk, MAX1LayerFinish, MAX1LayerStart
, Final_F1_0, Final_F1_1 , Final_F1_2 , Final_F1_3 , Final_F1_4 , Final_F1_5 , Final_F1_6 , Final_F1_7 , Final_F1_8 , Final_F1_9 , Final_F1_10 , Final_F1_11 , Final_F1_12 , Final_F1_13 , Final_F1_14 , Final_F1_15 , Final_F1_16 , Final_F1_17 , Final_F1_18 , Final_F1_19 , Final_F1_20 , Final_F1_21 , Final_F1_22 , Final_F1_23 , Final_F1_24 , Final_F1_25 , Final_F1_26 , Final_F1_27 , Final_F1_28 , Final_F1_29 , Final_F1_30 , Final_F1_31 , Final_F1_32 , Final_F1_33 , Final_F1_34 , Final_F1_35 , Final_F1_36 , Final_F1_37 , Final_F1_38 , Final_F1_39 , Final_F1_40 , Final_F1_41 , Final_F1_42 , Final_F1_43 , Final_F1_44 , Final_F1_45 , Final_F1_46 , Final_F1_47 , Final_F1_48 , Final_F1_49 , Final_F1_50 , Final_F1_51 , Final_F1_52 , Final_F1_53 , Final_F1_54 , Final_F1_55 , Final_F1_56 , Final_F1_57 , Final_F1_58 , Final_F1_59 , Final_F1_60 , Final_F1_61 , Final_F1_62 , Final_F1_63 , Final_F1_64 , Final_F1_65 , Final_F1_66 , Final_F1_67 , Final_F1_68 , Final_F1_69 , Final_F1_70 , Final_F1_71 , Final_F1_72 , Final_F1_73 , Final_F1_74 , Final_F1_75 , Final_F1_76 , Final_F1_77 , Final_F1_78 , Final_F1_79 , Final_F1_80 , Final_F1_81 , Final_F1_82 , Final_F1_83 , Final_F1_84 , Final_F1_85 , Final_F1_86 , Final_F1_87 , Final_F1_88 , Final_F1_89 , Final_F1_90 , Final_F1_91 , Final_F1_92 , Final_F1_93 , Final_F1_94 , Final_F1_95 , Final_F1_96 , Final_F1_97 , Final_F1_98 , Final_F1_99 , Final_F1_100 , Final_F1_101 , Final_F1_102 , Final_F1_103 , Final_F1_104 , Final_F1_105 , Final_F1_106 , Final_F1_107 , Final_F1_108 , Final_F1_109 , Final_F1_110 , Final_F1_111 , Final_F1_112 , Final_F1_113 , Final_F1_114 , Final_F1_115 , Final_F1_116 , Final_F1_117 , Final_F1_118 , Final_F1_119 , Final_F1_120 , Final_F1_121 , Final_F1_122 , Final_F1_123 , Final_F1_124 , Final_F1_125 , Final_F1_126 , Final_F1_127 , Final_F1_128 , Final_F1_129 , Final_F1_130 , Final_F1_131 , Final_F1_132 , Final_F1_133 , Final_F1_134 , Final_F1_135 , Final_F1_136 , Final_F1_137 , Final_F1_138 , Final_F1_139 , Final_F1_140 , Final_F1_141 , Final_F1_142 , Final_F1_143 , Final_F1_144 , Final_F1_145 , Final_F1_146 , Final_F1_147 , Final_F1_148 , Final_F1_149 , Final_F1_150 , Final_F1_151 , Final_F1_152 , Final_F1_153 , Final_F1_154 , Final_F1_155 , Final_F1_156 , Final_F1_157 , Final_F1_158 , Final_F1_159 , Final_F1_160 , Final_F1_161 , Final_F1_162 , Final_F1_163 , Final_F1_164 , Final_F1_165 , Final_F1_166 , Final_F1_167 , Final_F1_168 , Final_F1_169 , Final_F1_170 , Final_F1_171 , Final_F1_172 , Final_F1_173 , Final_F1_174 , Final_F1_175 , Final_F1_176 , Final_F1_177 , Final_F1_178 , Final_F1_179 , Final_F1_180 , Final_F1_181 , Final_F1_182 , Final_F1_183 , Final_F1_184 , Final_F1_185 , Final_F1_186 , Final_F1_187 , Final_F1_188 , Final_F1_189 , Final_F1_190 , Final_F1_191 , Final_F1_192 , Final_F1_193 , Final_F1_194 , Final_F1_195 , Final_F1_196 , Final_F1_197 , Final_F1_198 , Final_F1_199 , Final_F1_200 , Final_F1_201 , Final_F1_202 , Final_F1_203 , Final_F1_204 , Final_F1_205 , Final_F1_206 , Final_F1_207 , Final_F1_208 , Final_F1_209 , Final_F1_210 , Final_F1_211 , Final_F1_212 , Final_F1_213 , Final_F1_214 , Final_F1_215 , Final_F1_216 , Final_F1_217 , Final_F1_218 , Final_F1_219 , Final_F1_220 , Final_F1_221 , Final_F1_222 , Final_F1_223 , Final_F1_224 , Final_F1_225 , Final_F1_226 , Final_F1_227 , Final_F1_228 , Final_F1_229 , Final_F1_230 , Final_F1_231 , Final_F1_232 , Final_F1_233 , Final_F1_234 , Final_F1_235 , Final_F1_236 , Final_F1_237 , Final_F1_238 , Final_F1_239 , Final_F1_240 , Final_F1_241 , Final_F1_242 , Final_F1_243 , Final_F1_244 , Final_F1_245 , Final_F1_246 , Final_F1_247 , Final_F1_248 , Final_F1_249 , Final_F1_250 , Final_F1_251 , Final_F1_252 , Final_F1_253 , Final_F1_254 , Final_F1_255 , Final_F1_256 , Final_F1_257 , Final_F1_258 , Final_F1_259 , Final_F1_260 , Final_F1_261 , Final_F1_262 , Final_F1_263 , Final_F1_264 , Final_F1_265 , Final_F1_266 , Final_F1_267 , Final_F1_268 , Final_F1_269 , Final_F1_270 , Final_F1_271 , Final_F1_272 , Final_F1_273 , Final_F1_274 , Final_F1_275 , Final_F1_276 , Final_F1_277 , Final_F1_278 , Final_F1_279 , Final_F1_280 , Final_F1_281 , Final_F1_282 , Final_F1_283 , Final_F1_284 , Final_F1_285 , Final_F1_286 , Final_F1_287 , Final_F1_288 , Final_F1_289 , Final_F1_290 , Final_F1_291 , Final_F1_292 , Final_F1_293 , Final_F1_294 , Final_F1_295 , Final_F1_296 , Final_F1_297 , Final_F1_298 , Final_F1_299 , Final_F1_300 , Final_F1_301 , Final_F1_302 , Final_F1_303 , Final_F1_304 , Final_F1_305 , Final_F1_306 , Final_F1_307 , Final_F1_308 , Final_F1_309 , Final_F1_310 , Final_F1_311 , Final_F1_312 , Final_F1_313 , Final_F1_314 , Final_F1_315 , Final_F1_316 , Final_F1_317 , Final_F1_318 , Final_F1_319 , Final_F1_320 , Final_F1_321 , Final_F1_322 , Final_F1_323 , Final_F1_324 , Final_F1_325 , Final_F1_326 , Final_F1_327 , Final_F1_328 , Final_F1_329 , Final_F1_330 , Final_F1_331 , Final_F1_332 , Final_F1_333 , Final_F1_334 , Final_F1_335 , Final_F1_336 , Final_F1_337 , Final_F1_338 , Final_F1_339 , Final_F1_340 , Final_F1_341 , Final_F1_342 , Final_F1_343 , Final_F1_344 , Final_F1_345 , Final_F1_346 , Final_F1_347 , Final_F1_348 , Final_F1_349 , Final_F1_350 , Final_F1_351 , Final_F1_352 , Final_F1_353 , Final_F1_354 , Final_F1_355 , Final_F1_356 , Final_F1_357 , Final_F1_358 , Final_F1_359 , Final_F1_360 , Final_F1_361 , Final_F1_362 , Final_F1_363 , Final_F1_364 , Final_F1_365 , Final_F1_366 , Final_F1_367 , Final_F1_368 , Final_F1_369 , Final_F1_370 , Final_F1_371 , Final_F1_372 , Final_F1_373 , Final_F1_374 , Final_F1_375 , Final_F1_376 , Final_F1_377 , Final_F1_378 , Final_F1_379 , Final_F1_380 , Final_F1_381 , Final_F1_382 , Final_F1_383 , Final_F1_384 , Final_F1_385 , Final_F1_386 , Final_F1_387 , Final_F1_388 , Final_F1_389 , Final_F1_390 , Final_F1_391 , Final_F1_392 , Final_F1_393 , Final_F1_394 , Final_F1_395 , Final_F1_396 , Final_F1_397 , Final_F1_398 , Final_F1_399 , Final_F1_400 , Final_F1_401 , Final_F1_402 , Final_F1_403 , Final_F1_404 , Final_F1_405 , Final_F1_406 , Final_F1_407 , Final_F1_408 , Final_F1_409 , Final_F1_410 , Final_F1_411 , Final_F1_412 , Final_F1_413 , Final_F1_414 , Final_F1_415 , Final_F1_416 , Final_F1_417 , Final_F1_418 , Final_F1_419 , Final_F1_420 , Final_F1_421 , Final_F1_422 , Final_F1_423 , Final_F1_424 , Final_F1_425 , Final_F1_426 , Final_F1_427 , Final_F1_428 , Final_F1_429 , Final_F1_430 , Final_F1_431 , Final_F1_432 , Final_F1_433 , Final_F1_434 , Final_F1_435 , Final_F1_436 , Final_F1_437 , Final_F1_438 , Final_F1_439 , Final_F1_440 , Final_F1_441 , Final_F1_442 , Final_F1_443 , Final_F1_444 , Final_F1_445 , Final_F1_446 , Final_F1_447 , Final_F1_448 , Final_F1_449 , Final_F1_450 , Final_F1_451 , Final_F1_452 , Final_F1_453 , Final_F1_454 , Final_F1_455 , Final_F1_456 , Final_F1_457 , Final_F1_458 , Final_F1_459 , Final_F1_460 , Final_F1_461 , Final_F1_462 , Final_F1_463 , Final_F1_464 , Final_F1_465 , Final_F1_466 , Final_F1_467 , Final_F1_468 , Final_F1_469 , Final_F1_470 , Final_F1_471 , Final_F1_472 , Final_F1_473 , Final_F1_474 , Final_F1_475 , Final_F1_476 , Final_F1_477 , Final_F1_478 , Final_F1_479 , Final_F1_480 , Final_F1_481 , Final_F1_482 , Final_F1_483 , Final_F1_484 , Final_F1_485 , Final_F1_486 , Final_F1_487 , Final_F1_488 , Final_F1_489 , Final_F1_490 , Final_F1_491 , Final_F1_492 , Final_F1_493 , Final_F1_494 , Final_F1_495 , Final_F1_496 , Final_F1_497 , Final_F1_498 , Final_F1_499 , Final_F1_500 , Final_F1_501 , Final_F1_502 , Final_F1_503 , Final_F1_504 , Final_F1_505 , Final_F1_506 , Final_F1_507 , Final_F1_508 , Final_F1_509 , Final_F1_510 , Final_F1_511 , Final_F1_512 , Final_F1_513 , Final_F1_514 , Final_F1_515 , Final_F1_516 , Final_F1_517 , Final_F1_518 , Final_F1_519 , Final_F1_520 , Final_F1_521 , Final_F1_522 , Final_F1_523 , Final_F1_524 , Final_F1_525 , Final_F1_526 , Final_F1_527 , Final_F1_528 , Final_F1_529 , Final_F1_530 , Final_F1_531 , Final_F1_532 , Final_F1_533 , Final_F1_534 , Final_F1_535 , Final_F1_536 , Final_F1_537 , Final_F1_538 , Final_F1_539 , Final_F1_540 , Final_F1_541 , Final_F1_542 , Final_F1_543 , Final_F1_544 , Final_F1_545 , Final_F1_546 , Final_F1_547 , Final_F1_548 , Final_F1_549 , Final_F1_550 , Final_F1_551 , Final_F1_552 , Final_F1_553 , Final_F1_554 , Final_F1_555 , Final_F1_556 , Final_F1_557 , Final_F1_558 , Final_F1_559 , Final_F1_560 , Final_F1_561 , Final_F1_562 , Final_F1_563 , Final_F1_564 , Final_F1_565 , Final_F1_566 , Final_F1_567 , Final_F1_568 , Final_F1_569 , Final_F1_570 , Final_F1_571 , Final_F1_572 , Final_F1_573 , Final_F1_574 , Final_F1_575 
, Final_F2_0, Final_F2_1 , Final_F2_2 , Final_F2_3 , Final_F2_4 , Final_F2_5 , Final_F2_6 , Final_F2_7 , Final_F2_8 , Final_F2_9 , Final_F2_10 , Final_F2_11 , Final_F2_12 , Final_F2_13 , Final_F2_14 , Final_F2_15 , Final_F2_16 , Final_F2_17 , Final_F2_18 , Final_F2_19 , Final_F2_20 , Final_F2_21 , Final_F2_22 , Final_F2_23 , Final_F2_24 , Final_F2_25 , Final_F2_26 , Final_F2_27 , Final_F2_28 , Final_F2_29 , Final_F2_30 , Final_F2_31 , Final_F2_32 , Final_F2_33 , Final_F2_34 , Final_F2_35 , Final_F2_36 , Final_F2_37 , Final_F2_38 , Final_F2_39 , Final_F2_40 , Final_F2_41 , Final_F2_42 , Final_F2_43 , Final_F2_44 , Final_F2_45 , Final_F2_46 , Final_F2_47 , Final_F2_48 , Final_F2_49 , Final_F2_50 , Final_F2_51 , Final_F2_52 , Final_F2_53 , Final_F2_54 , Final_F2_55 , Final_F2_56 , Final_F2_57 , Final_F2_58 , Final_F2_59 , Final_F2_60 , Final_F2_61 , Final_F2_62 , Final_F2_63 , Final_F2_64 , Final_F2_65 , Final_F2_66 , Final_F2_67 , Final_F2_68 , Final_F2_69 , Final_F2_70 , Final_F2_71 , Final_F2_72 , Final_F2_73 , Final_F2_74 , Final_F2_75 , Final_F2_76 , Final_F2_77 , Final_F2_78 , Final_F2_79 , Final_F2_80 , Final_F2_81 , Final_F2_82 , Final_F2_83 , Final_F2_84 , Final_F2_85 , Final_F2_86 , Final_F2_87 , Final_F2_88 , Final_F2_89 , Final_F2_90 , Final_F2_91 , Final_F2_92 , Final_F2_93 , Final_F2_94 , Final_F2_95 , Final_F2_96 , Final_F2_97 , Final_F2_98 , Final_F2_99 , Final_F2_100 , Final_F2_101 , Final_F2_102 , Final_F2_103 , Final_F2_104 , Final_F2_105 , Final_F2_106 , Final_F2_107 , Final_F2_108 , Final_F2_109 , Final_F2_110 , Final_F2_111 , Final_F2_112 , Final_F2_113 , Final_F2_114 , Final_F2_115 , Final_F2_116 , Final_F2_117 , Final_F2_118 , Final_F2_119 , Final_F2_120 , Final_F2_121 , Final_F2_122 , Final_F2_123 , Final_F2_124 , Final_F2_125 , Final_F2_126 , Final_F2_127 , Final_F2_128 , Final_F2_129 , Final_F2_130 , Final_F2_131 , Final_F2_132 , Final_F2_133 , Final_F2_134 , Final_F2_135 , Final_F2_136 , Final_F2_137 , Final_F2_138 , Final_F2_139 , Final_F2_140 , Final_F2_141 , Final_F2_142 , Final_F2_143 , Final_F2_144 , Final_F2_145 , Final_F2_146 , Final_F2_147 , Final_F2_148 , Final_F2_149 , Final_F2_150 , Final_F2_151 , Final_F2_152 , Final_F2_153 , Final_F2_154 , Final_F2_155 , Final_F2_156 , Final_F2_157 , Final_F2_158 , Final_F2_159 , Final_F2_160 , Final_F2_161 , Final_F2_162 , Final_F2_163 , Final_F2_164 , Final_F2_165 , Final_F2_166 , Final_F2_167 , Final_F2_168 , Final_F2_169 , Final_F2_170 , Final_F2_171 , Final_F2_172 , Final_F2_173 , Final_F2_174 , Final_F2_175 , Final_F2_176 , Final_F2_177 , Final_F2_178 , Final_F2_179 , Final_F2_180 , Final_F2_181 , Final_F2_182 , Final_F2_183 , Final_F2_184 , Final_F2_185 , Final_F2_186 , Final_F2_187 , Final_F2_188 , Final_F2_189 , Final_F2_190 , Final_F2_191 , Final_F2_192 , Final_F2_193 , Final_F2_194 , Final_F2_195 , Final_F2_196 , Final_F2_197 , Final_F2_198 , Final_F2_199 , Final_F2_200 , Final_F2_201 , Final_F2_202 , Final_F2_203 , Final_F2_204 , Final_F2_205 , Final_F2_206 , Final_F2_207 , Final_F2_208 , Final_F2_209 , Final_F2_210 , Final_F2_211 , Final_F2_212 , Final_F2_213 , Final_F2_214 , Final_F2_215 , Final_F2_216 , Final_F2_217 , Final_F2_218 , Final_F2_219 , Final_F2_220 , Final_F2_221 , Final_F2_222 , Final_F2_223 , Final_F2_224 , Final_F2_225 , Final_F2_226 , Final_F2_227 , Final_F2_228 , Final_F2_229 , Final_F2_230 , Final_F2_231 , Final_F2_232 , Final_F2_233 , Final_F2_234 , Final_F2_235 , Final_F2_236 , Final_F2_237 , Final_F2_238 , Final_F2_239 , Final_F2_240 , Final_F2_241 , Final_F2_242 , Final_F2_243 , Final_F2_244 , Final_F2_245 , Final_F2_246 , Final_F2_247 , Final_F2_248 , Final_F2_249 , Final_F2_250 , Final_F2_251 , Final_F2_252 , Final_F2_253 , Final_F2_254 , Final_F2_255 , Final_F2_256 , Final_F2_257 , Final_F2_258 , Final_F2_259 , Final_F2_260 , Final_F2_261 , Final_F2_262 , Final_F2_263 , Final_F2_264 , Final_F2_265 , Final_F2_266 , Final_F2_267 , Final_F2_268 , Final_F2_269 , Final_F2_270 , Final_F2_271 , Final_F2_272 , Final_F2_273 , Final_F2_274 , Final_F2_275 , Final_F2_276 , Final_F2_277 , Final_F2_278 , Final_F2_279 , Final_F2_280 , Final_F2_281 , Final_F2_282 , Final_F2_283 , Final_F2_284 , Final_F2_285 , Final_F2_286 , Final_F2_287 , Final_F2_288 , Final_F2_289 , Final_F2_290 , Final_F2_291 , Final_F2_292 , Final_F2_293 , Final_F2_294 , Final_F2_295 , Final_F2_296 , Final_F2_297 , Final_F2_298 , Final_F2_299 , Final_F2_300 , Final_F2_301 , Final_F2_302 , Final_F2_303 , Final_F2_304 , Final_F2_305 , Final_F2_306 , Final_F2_307 , Final_F2_308 , Final_F2_309 , Final_F2_310 , Final_F2_311 , Final_F2_312 , Final_F2_313 , Final_F2_314 , Final_F2_315 , Final_F2_316 , Final_F2_317 , Final_F2_318 , Final_F2_319 , Final_F2_320 , Final_F2_321 , Final_F2_322 , Final_F2_323 , Final_F2_324 , Final_F2_325 , Final_F2_326 , Final_F2_327 , Final_F2_328 , Final_F2_329 , Final_F2_330 , Final_F2_331 , Final_F2_332 , Final_F2_333 , Final_F2_334 , Final_F2_335 , Final_F2_336 , Final_F2_337 , Final_F2_338 , Final_F2_339 , Final_F2_340 , Final_F2_341 , Final_F2_342 , Final_F2_343 , Final_F2_344 , Final_F2_345 , Final_F2_346 , Final_F2_347 , Final_F2_348 , Final_F2_349 , Final_F2_350 , Final_F2_351 , Final_F2_352 , Final_F2_353 , Final_F2_354 , Final_F2_355 , Final_F2_356 , Final_F2_357 , Final_F2_358 , Final_F2_359 , Final_F2_360 , Final_F2_361 , Final_F2_362 , Final_F2_363 , Final_F2_364 , Final_F2_365 , Final_F2_366 , Final_F2_367 , Final_F2_368 , Final_F2_369 , Final_F2_370 , Final_F2_371 , Final_F2_372 , Final_F2_373 , Final_F2_374 , Final_F2_375 , Final_F2_376 , Final_F2_377 , Final_F2_378 , Final_F2_379 , Final_F2_380 , Final_F2_381 , Final_F2_382 , Final_F2_383 , Final_F2_384 , Final_F2_385 , Final_F2_386 , Final_F2_387 , Final_F2_388 , Final_F2_389 , Final_F2_390 , Final_F2_391 , Final_F2_392 , Final_F2_393 , Final_F2_394 , Final_F2_395 , Final_F2_396 , Final_F2_397 , Final_F2_398 , Final_F2_399 , Final_F2_400 , Final_F2_401 , Final_F2_402 , Final_F2_403 , Final_F2_404 , Final_F2_405 , Final_F2_406 , Final_F2_407 , Final_F2_408 , Final_F2_409 , Final_F2_410 , Final_F2_411 , Final_F2_412 , Final_F2_413 , Final_F2_414 , Final_F2_415 , Final_F2_416 , Final_F2_417 , Final_F2_418 , Final_F2_419 , Final_F2_420 , Final_F2_421 , Final_F2_422 , Final_F2_423 , Final_F2_424 , Final_F2_425 , Final_F2_426 , Final_F2_427 , Final_F2_428 , Final_F2_429 , Final_F2_430 , Final_F2_431 , Final_F2_432 , Final_F2_433 , Final_F2_434 , Final_F2_435 , Final_F2_436 , Final_F2_437 , Final_F2_438 , Final_F2_439 , Final_F2_440 , Final_F2_441 , Final_F2_442 , Final_F2_443 , Final_F2_444 , Final_F2_445 , Final_F2_446 , Final_F2_447 , Final_F2_448 , Final_F2_449 , Final_F2_450 , Final_F2_451 , Final_F2_452 , Final_F2_453 , Final_F2_454 , Final_F2_455 , Final_F2_456 , Final_F2_457 , Final_F2_458 , Final_F2_459 , Final_F2_460 , Final_F2_461 , Final_F2_462 , Final_F2_463 , Final_F2_464 , Final_F2_465 , Final_F2_466 , Final_F2_467 , Final_F2_468 , Final_F2_469 , Final_F2_470 , Final_F2_471 , Final_F2_472 , Final_F2_473 , Final_F2_474 , Final_F2_475 , Final_F2_476 , Final_F2_477 , Final_F2_478 , Final_F2_479 , Final_F2_480 , Final_F2_481 , Final_F2_482 , Final_F2_483 , Final_F2_484 , Final_F2_485 , Final_F2_486 , Final_F2_487 , Final_F2_488 , Final_F2_489 , Final_F2_490 , Final_F2_491 , Final_F2_492 , Final_F2_493 , Final_F2_494 , Final_F2_495 , Final_F2_496 , Final_F2_497 , Final_F2_498 , Final_F2_499 , Final_F2_500 , Final_F2_501 , Final_F2_502 , Final_F2_503 , Final_F2_504 , Final_F2_505 , Final_F2_506 , Final_F2_507 , Final_F2_508 , Final_F2_509 , Final_F2_510 , Final_F2_511 , Final_F2_512 , Final_F2_513 , Final_F2_514 , Final_F2_515 , Final_F2_516 , Final_F2_517 , Final_F2_518 , Final_F2_519 , Final_F2_520 , Final_F2_521 , Final_F2_522 , Final_F2_523 , Final_F2_524 , Final_F2_525 , Final_F2_526 , Final_F2_527 , Final_F2_528 , Final_F2_529 , Final_F2_530 , Final_F2_531 , Final_F2_532 , Final_F2_533 , Final_F2_534 , Final_F2_535 , Final_F2_536 , Final_F2_537 , Final_F2_538 , Final_F2_539 , Final_F2_540 , Final_F2_541 , Final_F2_542 , Final_F2_543 , Final_F2_544 , Final_F2_545 , Final_F2_546 , Final_F2_547 , Final_F2_548 , Final_F2_549 , Final_F2_550 , Final_F2_551 , Final_F2_552 , Final_F2_553 , Final_F2_554 , Final_F2_555 , Final_F2_556 , Final_F2_557 , Final_F2_558 , Final_F2_559 , Final_F2_560 , Final_F2_561 , Final_F2_562 , Final_F2_563 , Final_F2_564 , Final_F2_565 , Final_F2_566 , Final_F2_567 , Final_F2_568 , Final_F2_569 , Final_F2_570 , Final_F2_571 , Final_F2_572 , Final_F2_573 , Final_F2_574 , Final_F2_575 
, Final_F3_0, Final_F3_1 , Final_F3_2 , Final_F3_3 , Final_F3_4 , Final_F3_5 , Final_F3_6 , Final_F3_7 , Final_F3_8 , Final_F3_9 , Final_F3_10 , Final_F3_11 , Final_F3_12 , Final_F3_13 , Final_F3_14 , Final_F3_15 , Final_F3_16 , Final_F3_17 , Final_F3_18 , Final_F3_19 , Final_F3_20 , Final_F3_21 , Final_F3_22 , Final_F3_23 , Final_F3_24 , Final_F3_25 , Final_F3_26 , Final_F3_27 , Final_F3_28 , Final_F3_29 , Final_F3_30 , Final_F3_31 , Final_F3_32 , Final_F3_33 , Final_F3_34 , Final_F3_35 , Final_F3_36 , Final_F3_37 , Final_F3_38 , Final_F3_39 , Final_F3_40 , Final_F3_41 , Final_F3_42 , Final_F3_43 , Final_F3_44 , Final_F3_45 , Final_F3_46 , Final_F3_47 , Final_F3_48 , Final_F3_49 , Final_F3_50 , Final_F3_51 , Final_F3_52 , Final_F3_53 , Final_F3_54 , Final_F3_55 , Final_F3_56 , Final_F3_57 , Final_F3_58 , Final_F3_59 , Final_F3_60 , Final_F3_61 , Final_F3_62 , Final_F3_63 , Final_F3_64 , Final_F3_65 , Final_F3_66 , Final_F3_67 , Final_F3_68 , Final_F3_69 , Final_F3_70 , Final_F3_71 , Final_F3_72 , Final_F3_73 , Final_F3_74 , Final_F3_75 , Final_F3_76 , Final_F3_77 , Final_F3_78 , Final_F3_79 , Final_F3_80 , Final_F3_81 , Final_F3_82 , Final_F3_83 , Final_F3_84 , Final_F3_85 , Final_F3_86 , Final_F3_87 , Final_F3_88 , Final_F3_89 , Final_F3_90 , Final_F3_91 , Final_F3_92 , Final_F3_93 , Final_F3_94 , Final_F3_95 , Final_F3_96 , Final_F3_97 , Final_F3_98 , Final_F3_99 , Final_F3_100 , Final_F3_101 , Final_F3_102 , Final_F3_103 , Final_F3_104 , Final_F3_105 , Final_F3_106 , Final_F3_107 , Final_F3_108 , Final_F3_109 , Final_F3_110 , Final_F3_111 , Final_F3_112 , Final_F3_113 , Final_F3_114 , Final_F3_115 , Final_F3_116 , Final_F3_117 , Final_F3_118 , Final_F3_119 , Final_F3_120 , Final_F3_121 , Final_F3_122 , Final_F3_123 , Final_F3_124 , Final_F3_125 , Final_F3_126 , Final_F3_127 , Final_F3_128 , Final_F3_129 , Final_F3_130 , Final_F3_131 , Final_F3_132 , Final_F3_133 , Final_F3_134 , Final_F3_135 , Final_F3_136 , Final_F3_137 , Final_F3_138 , Final_F3_139 , Final_F3_140 , Final_F3_141 , Final_F3_142 , Final_F3_143 , Final_F3_144 , Final_F3_145 , Final_F3_146 , Final_F3_147 , Final_F3_148 , Final_F3_149 , Final_F3_150 , Final_F3_151 , Final_F3_152 , Final_F3_153 , Final_F3_154 , Final_F3_155 , Final_F3_156 , Final_F3_157 , Final_F3_158 , Final_F3_159 , Final_F3_160 , Final_F3_161 , Final_F3_162 , Final_F3_163 , Final_F3_164 , Final_F3_165 , Final_F3_166 , Final_F3_167 , Final_F3_168 , Final_F3_169 , Final_F3_170 , Final_F3_171 , Final_F3_172 , Final_F3_173 , Final_F3_174 , Final_F3_175 , Final_F3_176 , Final_F3_177 , Final_F3_178 , Final_F3_179 , Final_F3_180 , Final_F3_181 , Final_F3_182 , Final_F3_183 , Final_F3_184 , Final_F3_185 , Final_F3_186 , Final_F3_187 , Final_F3_188 , Final_F3_189 , Final_F3_190 , Final_F3_191 , Final_F3_192 , Final_F3_193 , Final_F3_194 , Final_F3_195 , Final_F3_196 , Final_F3_197 , Final_F3_198 , Final_F3_199 , Final_F3_200 , Final_F3_201 , Final_F3_202 , Final_F3_203 , Final_F3_204 , Final_F3_205 , Final_F3_206 , Final_F3_207 , Final_F3_208 , Final_F3_209 , Final_F3_210 , Final_F3_211 , Final_F3_212 , Final_F3_213 , Final_F3_214 , Final_F3_215 , Final_F3_216 , Final_F3_217 , Final_F3_218 , Final_F3_219 , Final_F3_220 , Final_F3_221 , Final_F3_222 , Final_F3_223 , Final_F3_224 , Final_F3_225 , Final_F3_226 , Final_F3_227 , Final_F3_228 , Final_F3_229 , Final_F3_230 , Final_F3_231 , Final_F3_232 , Final_F3_233 , Final_F3_234 , Final_F3_235 , Final_F3_236 , Final_F3_237 , Final_F3_238 , Final_F3_239 , Final_F3_240 , Final_F3_241 , Final_F3_242 , Final_F3_243 , Final_F3_244 , Final_F3_245 , Final_F3_246 , Final_F3_247 , Final_F3_248 , Final_F3_249 , Final_F3_250 , Final_F3_251 , Final_F3_252 , Final_F3_253 , Final_F3_254 , Final_F3_255 , Final_F3_256 , Final_F3_257 , Final_F3_258 , Final_F3_259 , Final_F3_260 , Final_F3_261 , Final_F3_262 , Final_F3_263 , Final_F3_264 , Final_F3_265 , Final_F3_266 , Final_F3_267 , Final_F3_268 , Final_F3_269 , Final_F3_270 , Final_F3_271 , Final_F3_272 , Final_F3_273 , Final_F3_274 , Final_F3_275 , Final_F3_276 , Final_F3_277 , Final_F3_278 , Final_F3_279 , Final_F3_280 , Final_F3_281 , Final_F3_282 , Final_F3_283 , Final_F3_284 , Final_F3_285 , Final_F3_286 , Final_F3_287 , Final_F3_288 , Final_F3_289 , Final_F3_290 , Final_F3_291 , Final_F3_292 , Final_F3_293 , Final_F3_294 , Final_F3_295 , Final_F3_296 , Final_F3_297 , Final_F3_298 , Final_F3_299 , Final_F3_300 , Final_F3_301 , Final_F3_302 , Final_F3_303 , Final_F3_304 , Final_F3_305 , Final_F3_306 , Final_F3_307 , Final_F3_308 , Final_F3_309 , Final_F3_310 , Final_F3_311 , Final_F3_312 , Final_F3_313 , Final_F3_314 , Final_F3_315 , Final_F3_316 , Final_F3_317 , Final_F3_318 , Final_F3_319 , Final_F3_320 , Final_F3_321 , Final_F3_322 , Final_F3_323 , Final_F3_324 , Final_F3_325 , Final_F3_326 , Final_F3_327 , Final_F3_328 , Final_F3_329 , Final_F3_330 , Final_F3_331 , Final_F3_332 , Final_F3_333 , Final_F3_334 , Final_F3_335 , Final_F3_336 , Final_F3_337 , Final_F3_338 , Final_F3_339 , Final_F3_340 , Final_F3_341 , Final_F3_342 , Final_F3_343 , Final_F3_344 , Final_F3_345 , Final_F3_346 , Final_F3_347 , Final_F3_348 , Final_F3_349 , Final_F3_350 , Final_F3_351 , Final_F3_352 , Final_F3_353 , Final_F3_354 , Final_F3_355 , Final_F3_356 , Final_F3_357 , Final_F3_358 , Final_F3_359 , Final_F3_360 , Final_F3_361 , Final_F3_362 , Final_F3_363 , Final_F3_364 , Final_F3_365 , Final_F3_366 , Final_F3_367 , Final_F3_368 , Final_F3_369 , Final_F3_370 , Final_F3_371 , Final_F3_372 , Final_F3_373 , Final_F3_374 , Final_F3_375 , Final_F3_376 , Final_F3_377 , Final_F3_378 , Final_F3_379 , Final_F3_380 , Final_F3_381 , Final_F3_382 , Final_F3_383 , Final_F3_384 , Final_F3_385 , Final_F3_386 , Final_F3_387 , Final_F3_388 , Final_F3_389 , Final_F3_390 , Final_F3_391 , Final_F3_392 , Final_F3_393 , Final_F3_394 , Final_F3_395 , Final_F3_396 , Final_F3_397 , Final_F3_398 , Final_F3_399 , Final_F3_400 , Final_F3_401 , Final_F3_402 , Final_F3_403 , Final_F3_404 , Final_F3_405 , Final_F3_406 , Final_F3_407 , Final_F3_408 , Final_F3_409 , Final_F3_410 , Final_F3_411 , Final_F3_412 , Final_F3_413 , Final_F3_414 , Final_F3_415 , Final_F3_416 , Final_F3_417 , Final_F3_418 , Final_F3_419 , Final_F3_420 , Final_F3_421 , Final_F3_422 , Final_F3_423 , Final_F3_424 , Final_F3_425 , Final_F3_426 , Final_F3_427 , Final_F3_428 , Final_F3_429 , Final_F3_430 , Final_F3_431 , Final_F3_432 , Final_F3_433 , Final_F3_434 , Final_F3_435 , Final_F3_436 , Final_F3_437 , Final_F3_438 , Final_F3_439 , Final_F3_440 , Final_F3_441 , Final_F3_442 , Final_F3_443 , Final_F3_444 , Final_F3_445 , Final_F3_446 , Final_F3_447 , Final_F3_448 , Final_F3_449 , Final_F3_450 , Final_F3_451 , Final_F3_452 , Final_F3_453 , Final_F3_454 , Final_F3_455 , Final_F3_456 , Final_F3_457 , Final_F3_458 , Final_F3_459 , Final_F3_460 , Final_F3_461 , Final_F3_462 , Final_F3_463 , Final_F3_464 , Final_F3_465 , Final_F3_466 , Final_F3_467 , Final_F3_468 , Final_F3_469 , Final_F3_470 , Final_F3_471 , Final_F3_472 , Final_F3_473 , Final_F3_474 , Final_F3_475 , Final_F3_476 , Final_F3_477 , Final_F3_478 , Final_F3_479 , Final_F3_480 , Final_F3_481 , Final_F3_482 , Final_F3_483 , Final_F3_484 , Final_F3_485 , Final_F3_486 , Final_F3_487 , Final_F3_488 , Final_F3_489 , Final_F3_490 , Final_F3_491 , Final_F3_492 , Final_F3_493 , Final_F3_494 , Final_F3_495 , Final_F3_496 , Final_F3_497 , Final_F3_498 , Final_F3_499 , Final_F3_500 , Final_F3_501 , Final_F3_502 , Final_F3_503 , Final_F3_504 , Final_F3_505 , Final_F3_506 , Final_F3_507 , Final_F3_508 , Final_F3_509 , Final_F3_510 , Final_F3_511 , Final_F3_512 , Final_F3_513 , Final_F3_514 , Final_F3_515 , Final_F3_516 , Final_F3_517 , Final_F3_518 , Final_F3_519 , Final_F3_520 , Final_F3_521 , Final_F3_522 , Final_F3_523 , Final_F3_524 , Final_F3_525 , Final_F3_526 , Final_F3_527 , Final_F3_528 , Final_F3_529 , Final_F3_530 , Final_F3_531 , Final_F3_532 , Final_F3_533 , Final_F3_534 , Final_F3_535 , Final_F3_536 , Final_F3_537 , Final_F3_538 , Final_F3_539 , Final_F3_540 , Final_F3_541 , Final_F3_542 , Final_F3_543 , Final_F3_544 , Final_F3_545 , Final_F3_546 , Final_F3_547 , Final_F3_548 , Final_F3_549 , Final_F3_550 , Final_F3_551 , Final_F3_552 , Final_F3_553 , Final_F3_554 , Final_F3_555 , Final_F3_556 , Final_F3_557 , Final_F3_558 , Final_F3_559 , Final_F3_560 , Final_F3_561 , Final_F3_562 , Final_F3_563 , Final_F3_564 , Final_F3_565 , Final_F3_566 , Final_F3_567 , Final_F3_568 , Final_F3_569 , Final_F3_570 , Final_F3_571 , Final_F3_572 , Final_F3_573 , Final_F3_574 , Final_F3_575 
, Final_F4_0, Final_F4_1 , Final_F4_2 , Final_F4_3 , Final_F4_4 , Final_F4_5 , Final_F4_6 , Final_F4_7 , Final_F4_8 , Final_F4_9 , Final_F4_10 , Final_F4_11 , Final_F4_12 , Final_F4_13 , Final_F4_14 , Final_F4_15 , Final_F4_16 , Final_F4_17 , Final_F4_18 , Final_F4_19 , Final_F4_20 , Final_F4_21 , Final_F4_22 , Final_F4_23 , Final_F4_24 , Final_F4_25 , Final_F4_26 , Final_F4_27 , Final_F4_28 , Final_F4_29 , Final_F4_30 , Final_F4_31 , Final_F4_32 , Final_F4_33 , Final_F4_34 , Final_F4_35 , Final_F4_36 , Final_F4_37 , Final_F4_38 , Final_F4_39 , Final_F4_40 , Final_F4_41 , Final_F4_42 , Final_F4_43 , Final_F4_44 , Final_F4_45 , Final_F4_46 , Final_F4_47 , Final_F4_48 , Final_F4_49 , Final_F4_50 , Final_F4_51 , Final_F4_52 , Final_F4_53 , Final_F4_54 , Final_F4_55 , Final_F4_56 , Final_F4_57 , Final_F4_58 , Final_F4_59 , Final_F4_60 , Final_F4_61 , Final_F4_62 , Final_F4_63 , Final_F4_64 , Final_F4_65 , Final_F4_66 , Final_F4_67 , Final_F4_68 , Final_F4_69 , Final_F4_70 , Final_F4_71 , Final_F4_72 , Final_F4_73 , Final_F4_74 , Final_F4_75 , Final_F4_76 , Final_F4_77 , Final_F4_78 , Final_F4_79 , Final_F4_80 , Final_F4_81 , Final_F4_82 , Final_F4_83 , Final_F4_84 , Final_F4_85 , Final_F4_86 , Final_F4_87 , Final_F4_88 , Final_F4_89 , Final_F4_90 , Final_F4_91 , Final_F4_92 , Final_F4_93 , Final_F4_94 , Final_F4_95 , Final_F4_96 , Final_F4_97 , Final_F4_98 , Final_F4_99 , Final_F4_100 , Final_F4_101 , Final_F4_102 , Final_F4_103 , Final_F4_104 , Final_F4_105 , Final_F4_106 , Final_F4_107 , Final_F4_108 , Final_F4_109 , Final_F4_110 , Final_F4_111 , Final_F4_112 , Final_F4_113 , Final_F4_114 , Final_F4_115 , Final_F4_116 , Final_F4_117 , Final_F4_118 , Final_F4_119 , Final_F4_120 , Final_F4_121 , Final_F4_122 , Final_F4_123 , Final_F4_124 , Final_F4_125 , Final_F4_126 , Final_F4_127 , Final_F4_128 , Final_F4_129 , Final_F4_130 , Final_F4_131 , Final_F4_132 , Final_F4_133 , Final_F4_134 , Final_F4_135 , Final_F4_136 , Final_F4_137 , Final_F4_138 , Final_F4_139 , Final_F4_140 , Final_F4_141 , Final_F4_142 , Final_F4_143 , Final_F4_144 , Final_F4_145 , Final_F4_146 , Final_F4_147 , Final_F4_148 , Final_F4_149 , Final_F4_150 , Final_F4_151 , Final_F4_152 , Final_F4_153 , Final_F4_154 , Final_F4_155 , Final_F4_156 , Final_F4_157 , Final_F4_158 , Final_F4_159 , Final_F4_160 , Final_F4_161 , Final_F4_162 , Final_F4_163 , Final_F4_164 , Final_F4_165 , Final_F4_166 , Final_F4_167 , Final_F4_168 , Final_F4_169 , Final_F4_170 , Final_F4_171 , Final_F4_172 , Final_F4_173 , Final_F4_174 , Final_F4_175 , Final_F4_176 , Final_F4_177 , Final_F4_178 , Final_F4_179 , Final_F4_180 , Final_F4_181 , Final_F4_182 , Final_F4_183 , Final_F4_184 , Final_F4_185 , Final_F4_186 , Final_F4_187 , Final_F4_188 , Final_F4_189 , Final_F4_190 , Final_F4_191 , Final_F4_192 , Final_F4_193 , Final_F4_194 , Final_F4_195 , Final_F4_196 , Final_F4_197 , Final_F4_198 , Final_F4_199 , Final_F4_200 , Final_F4_201 , Final_F4_202 , Final_F4_203 , Final_F4_204 , Final_F4_205 , Final_F4_206 , Final_F4_207 , Final_F4_208 , Final_F4_209 , Final_F4_210 , Final_F4_211 , Final_F4_212 , Final_F4_213 , Final_F4_214 , Final_F4_215 , Final_F4_216 , Final_F4_217 , Final_F4_218 , Final_F4_219 , Final_F4_220 , Final_F4_221 , Final_F4_222 , Final_F4_223 , Final_F4_224 , Final_F4_225 , Final_F4_226 , Final_F4_227 , Final_F4_228 , Final_F4_229 , Final_F4_230 , Final_F4_231 , Final_F4_232 , Final_F4_233 , Final_F4_234 , Final_F4_235 , Final_F4_236 , Final_F4_237 , Final_F4_238 , Final_F4_239 , Final_F4_240 , Final_F4_241 , Final_F4_242 , Final_F4_243 , Final_F4_244 , Final_F4_245 , Final_F4_246 , Final_F4_247 , Final_F4_248 , Final_F4_249 , Final_F4_250 , Final_F4_251 , Final_F4_252 , Final_F4_253 , Final_F4_254 , Final_F4_255 , Final_F4_256 , Final_F4_257 , Final_F4_258 , Final_F4_259 , Final_F4_260 , Final_F4_261 , Final_F4_262 , Final_F4_263 , Final_F4_264 , Final_F4_265 , Final_F4_266 , Final_F4_267 , Final_F4_268 , Final_F4_269 , Final_F4_270 , Final_F4_271 , Final_F4_272 , Final_F4_273 , Final_F4_274 , Final_F4_275 , Final_F4_276 , Final_F4_277 , Final_F4_278 , Final_F4_279 , Final_F4_280 , Final_F4_281 , Final_F4_282 , Final_F4_283 , Final_F4_284 , Final_F4_285 , Final_F4_286 , Final_F4_287 , Final_F4_288 , Final_F4_289 , Final_F4_290 , Final_F4_291 , Final_F4_292 , Final_F4_293 , Final_F4_294 , Final_F4_295 , Final_F4_296 , Final_F4_297 , Final_F4_298 , Final_F4_299 , Final_F4_300 , Final_F4_301 , Final_F4_302 , Final_F4_303 , Final_F4_304 , Final_F4_305 , Final_F4_306 , Final_F4_307 , Final_F4_308 , Final_F4_309 , Final_F4_310 , Final_F4_311 , Final_F4_312 , Final_F4_313 , Final_F4_314 , Final_F4_315 , Final_F4_316 , Final_F4_317 , Final_F4_318 , Final_F4_319 , Final_F4_320 , Final_F4_321 , Final_F4_322 , Final_F4_323 , Final_F4_324 , Final_F4_325 , Final_F4_326 , Final_F4_327 , Final_F4_328 , Final_F4_329 , Final_F4_330 , Final_F4_331 , Final_F4_332 , Final_F4_333 , Final_F4_334 , Final_F4_335 , Final_F4_336 , Final_F4_337 , Final_F4_338 , Final_F4_339 , Final_F4_340 , Final_F4_341 , Final_F4_342 , Final_F4_343 , Final_F4_344 , Final_F4_345 , Final_F4_346 , Final_F4_347 , Final_F4_348 , Final_F4_349 , Final_F4_350 , Final_F4_351 , Final_F4_352 , Final_F4_353 , Final_F4_354 , Final_F4_355 , Final_F4_356 , Final_F4_357 , Final_F4_358 , Final_F4_359 , Final_F4_360 , Final_F4_361 , Final_F4_362 , Final_F4_363 , Final_F4_364 , Final_F4_365 , Final_F4_366 , Final_F4_367 , Final_F4_368 , Final_F4_369 , Final_F4_370 , Final_F4_371 , Final_F4_372 , Final_F4_373 , Final_F4_374 , Final_F4_375 , Final_F4_376 , Final_F4_377 , Final_F4_378 , Final_F4_379 , Final_F4_380 , Final_F4_381 , Final_F4_382 , Final_F4_383 , Final_F4_384 , Final_F4_385 , Final_F4_386 , Final_F4_387 , Final_F4_388 , Final_F4_389 , Final_F4_390 , Final_F4_391 , Final_F4_392 , Final_F4_393 , Final_F4_394 , Final_F4_395 , Final_F4_396 , Final_F4_397 , Final_F4_398 , Final_F4_399 , Final_F4_400 , Final_F4_401 , Final_F4_402 , Final_F4_403 , Final_F4_404 , Final_F4_405 , Final_F4_406 , Final_F4_407 , Final_F4_408 , Final_F4_409 , Final_F4_410 , Final_F4_411 , Final_F4_412 , Final_F4_413 , Final_F4_414 , Final_F4_415 , Final_F4_416 , Final_F4_417 , Final_F4_418 , Final_F4_419 , Final_F4_420 , Final_F4_421 , Final_F4_422 , Final_F4_423 , Final_F4_424 , Final_F4_425 , Final_F4_426 , Final_F4_427 , Final_F4_428 , Final_F4_429 , Final_F4_430 , Final_F4_431 , Final_F4_432 , Final_F4_433 , Final_F4_434 , Final_F4_435 , Final_F4_436 , Final_F4_437 , Final_F4_438 , Final_F4_439 , Final_F4_440 , Final_F4_441 , Final_F4_442 , Final_F4_443 , Final_F4_444 , Final_F4_445 , Final_F4_446 , Final_F4_447 , Final_F4_448 , Final_F4_449 , Final_F4_450 , Final_F4_451 , Final_F4_452 , Final_F4_453 , Final_F4_454 , Final_F4_455 , Final_F4_456 , Final_F4_457 , Final_F4_458 , Final_F4_459 , Final_F4_460 , Final_F4_461 , Final_F4_462 , Final_F4_463 , Final_F4_464 , Final_F4_465 , Final_F4_466 , Final_F4_467 , Final_F4_468 , Final_F4_469 , Final_F4_470 , Final_F4_471 , Final_F4_472 , Final_F4_473 , Final_F4_474 , Final_F4_475 , Final_F4_476 , Final_F4_477 , Final_F4_478 , Final_F4_479 , Final_F4_480 , Final_F4_481 , Final_F4_482 , Final_F4_483 , Final_F4_484 , Final_F4_485 , Final_F4_486 , Final_F4_487 , Final_F4_488 , Final_F4_489 , Final_F4_490 , Final_F4_491 , Final_F4_492 , Final_F4_493 , Final_F4_494 , Final_F4_495 , Final_F4_496 , Final_F4_497 , Final_F4_498 , Final_F4_499 , Final_F4_500 , Final_F4_501 , Final_F4_502 , Final_F4_503 , Final_F4_504 , Final_F4_505 , Final_F4_506 , Final_F4_507 , Final_F4_508 , Final_F4_509 , Final_F4_510 , Final_F4_511 , Final_F4_512 , Final_F4_513 , Final_F4_514 , Final_F4_515 , Final_F4_516 , Final_F4_517 , Final_F4_518 , Final_F4_519 , Final_F4_520 , Final_F4_521 , Final_F4_522 , Final_F4_523 , Final_F4_524 , Final_F4_525 , Final_F4_526 , Final_F4_527 , Final_F4_528 , Final_F4_529 , Final_F4_530 , Final_F4_531 , Final_F4_532 , Final_F4_533 , Final_F4_534 , Final_F4_535 , Final_F4_536 , Final_F4_537 , Final_F4_538 , Final_F4_539 , Final_F4_540 , Final_F4_541 , Final_F4_542 , Final_F4_543 , Final_F4_544 , Final_F4_545 , Final_F4_546 , Final_F4_547 , Final_F4_548 , Final_F4_549 , Final_F4_550 , Final_F4_551 , Final_F4_552 , Final_F4_553 , Final_F4_554 , Final_F4_555 , Final_F4_556 , Final_F4_557 , Final_F4_558 , Final_F4_559 , Final_F4_560 , Final_F4_561 , Final_F4_562 , Final_F4_563 , Final_F4_564 , Final_F4_565 , Final_F4_566 , Final_F4_567 , Final_F4_568 , Final_F4_569 , Final_F4_570 , Final_F4_571 , Final_F4_572 , Final_F4_573 , Final_F4_574 , Final_F4_575 
,REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143 
);
 
input clk;
input MAX1LayerStart;
*/
//output MAX1LayerFinish;


/* wire[8:0]  superADDRESS;  */
/* 
input wire [65:0] Final_F1_0, Final_F1_1 , Final_F1_2 , Final_F1_3 , Final_F1_4 , Final_F1_5 , Final_F1_6 , Final_F1_7 , Final_F1_8 , Final_F1_9 , Final_F1_10 , Final_F1_11 , Final_F1_12 , Final_F1_13 , Final_F1_14 , Final_F1_15 , Final_F1_16 , Final_F1_17 , Final_F1_18 , Final_F1_19 , Final_F1_20 , Final_F1_21 , Final_F1_22 , Final_F1_23 , Final_F1_24 , Final_F1_25 , Final_F1_26 , Final_F1_27 , Final_F1_28 , Final_F1_29 , Final_F1_30 , Final_F1_31 , Final_F1_32 , Final_F1_33 , Final_F1_34 , Final_F1_35 , Final_F1_36 , Final_F1_37 , Final_F1_38 , Final_F1_39 , Final_F1_40 , Final_F1_41 , Final_F1_42 , Final_F1_43 , Final_F1_44 , Final_F1_45 , Final_F1_46 , Final_F1_47 , Final_F1_48 , Final_F1_49 , Final_F1_50 , Final_F1_51 , Final_F1_52 , Final_F1_53 , Final_F1_54 , Final_F1_55 , Final_F1_56 , Final_F1_57 , Final_F1_58 , Final_F1_59 , Final_F1_60 , Final_F1_61 , Final_F1_62 , Final_F1_63 , Final_F1_64 , Final_F1_65 , Final_F1_66 , Final_F1_67 , Final_F1_68 , Final_F1_69 , Final_F1_70 , Final_F1_71 , Final_F1_72 , Final_F1_73 , Final_F1_74 , Final_F1_75 , Final_F1_76 , Final_F1_77 , Final_F1_78 , Final_F1_79 , Final_F1_80 , Final_F1_81 , Final_F1_82 , Final_F1_83 , Final_F1_84 , Final_F1_85 , Final_F1_86 , Final_F1_87 , Final_F1_88 , Final_F1_89 , Final_F1_90 , Final_F1_91 , Final_F1_92 , Final_F1_93 , Final_F1_94 , Final_F1_95 , Final_F1_96 , Final_F1_97 , Final_F1_98 , Final_F1_99 , Final_F1_100 , Final_F1_101 , Final_F1_102 , Final_F1_103 , Final_F1_104 , Final_F1_105 , Final_F1_106 , Final_F1_107 , Final_F1_108 , Final_F1_109 , Final_F1_110 , Final_F1_111 , Final_F1_112 , Final_F1_113 , Final_F1_114 , Final_F1_115 , Final_F1_116 , Final_F1_117 , Final_F1_118 , Final_F1_119 , Final_F1_120 , Final_F1_121 , Final_F1_122 , Final_F1_123 , Final_F1_124 , Final_F1_125 , Final_F1_126 , Final_F1_127 , Final_F1_128 , Final_F1_129 , Final_F1_130 , Final_F1_131 , Final_F1_132 , Final_F1_133 , Final_F1_134 , Final_F1_135 , Final_F1_136 , Final_F1_137 , Final_F1_138 , Final_F1_139 , Final_F1_140 , Final_F1_141 , Final_F1_142 , Final_F1_143 , Final_F1_144 , Final_F1_145 , Final_F1_146 , Final_F1_147 , Final_F1_148 , Final_F1_149 , Final_F1_150 , Final_F1_151 , Final_F1_152 , Final_F1_153 , Final_F1_154 , Final_F1_155 , Final_F1_156 , Final_F1_157 , Final_F1_158 , Final_F1_159 , Final_F1_160 , Final_F1_161 , Final_F1_162 , Final_F1_163 , Final_F1_164 , Final_F1_165 , Final_F1_166 , Final_F1_167 , Final_F1_168 , Final_F1_169 , Final_F1_170 , Final_F1_171 , Final_F1_172 , Final_F1_173 , Final_F1_174 , Final_F1_175 , Final_F1_176 , Final_F1_177 , Final_F1_178 , Final_F1_179 , Final_F1_180 , Final_F1_181 , Final_F1_182 , Final_F1_183 , Final_F1_184 , Final_F1_185 , Final_F1_186 , Final_F1_187 , Final_F1_188 , Final_F1_189 , Final_F1_190 , Final_F1_191 , Final_F1_192 , Final_F1_193 , Final_F1_194 , Final_F1_195 , Final_F1_196 , Final_F1_197 , Final_F1_198 , Final_F1_199 , Final_F1_200 , Final_F1_201 , Final_F1_202 , Final_F1_203 , Final_F1_204 , Final_F1_205 , Final_F1_206 , Final_F1_207 , Final_F1_208 , Final_F1_209 , Final_F1_210 , Final_F1_211 , Final_F1_212 , Final_F1_213 , Final_F1_214 , Final_F1_215 , Final_F1_216 , Final_F1_217 , Final_F1_218 , Final_F1_219 , Final_F1_220 , Final_F1_221 , Final_F1_222 , Final_F1_223 , Final_F1_224 , Final_F1_225 , Final_F1_226 , Final_F1_227 , Final_F1_228 , Final_F1_229 , Final_F1_230 , Final_F1_231 , Final_F1_232 , Final_F1_233 , Final_F1_234 , Final_F1_235 , Final_F1_236 , Final_F1_237 , Final_F1_238 , Final_F1_239 , Final_F1_240 , Final_F1_241 , Final_F1_242 , Final_F1_243 , Final_F1_244 , Final_F1_245 , Final_F1_246 , Final_F1_247 , Final_F1_248 , Final_F1_249 , Final_F1_250 , Final_F1_251 , Final_F1_252 , Final_F1_253 , Final_F1_254 , Final_F1_255 , Final_F1_256 , Final_F1_257 , Final_F1_258 , Final_F1_259 , Final_F1_260 , Final_F1_261 , Final_F1_262 , Final_F1_263 , Final_F1_264 , Final_F1_265 , Final_F1_266 , Final_F1_267 , Final_F1_268 , Final_F1_269 , Final_F1_270 , Final_F1_271 , Final_F1_272 , Final_F1_273 , Final_F1_274 , Final_F1_275 , Final_F1_276 , Final_F1_277 , Final_F1_278 , Final_F1_279 , Final_F1_280 , Final_F1_281 , Final_F1_282 , Final_F1_283 , Final_F1_284 , Final_F1_285 , Final_F1_286 , Final_F1_287 , Final_F1_288 , Final_F1_289 , Final_F1_290 , Final_F1_291 , Final_F1_292 , Final_F1_293 , Final_F1_294 , Final_F1_295 , Final_F1_296 , Final_F1_297 , Final_F1_298 , Final_F1_299 , Final_F1_300 , Final_F1_301 , Final_F1_302 , Final_F1_303 , Final_F1_304 , Final_F1_305 , Final_F1_306 , Final_F1_307 , Final_F1_308 , Final_F1_309 , Final_F1_310 , Final_F1_311 , Final_F1_312 , Final_F1_313 , Final_F1_314 , Final_F1_315 , Final_F1_316 , Final_F1_317 , Final_F1_318 , Final_F1_319 , Final_F1_320 , Final_F1_321 , Final_F1_322 , Final_F1_323 , Final_F1_324 , Final_F1_325 , Final_F1_326 , Final_F1_327 , Final_F1_328 , Final_F1_329 , Final_F1_330 , Final_F1_331 , Final_F1_332 , Final_F1_333 , Final_F1_334 , Final_F1_335 , Final_F1_336 , Final_F1_337 , Final_F1_338 , Final_F1_339 , Final_F1_340 , Final_F1_341 , Final_F1_342 , Final_F1_343 , Final_F1_344 , Final_F1_345 , Final_F1_346 , Final_F1_347 , Final_F1_348 , Final_F1_349 , Final_F1_350 , Final_F1_351 , Final_F1_352 , Final_F1_353 , Final_F1_354 , Final_F1_355 , Final_F1_356 , Final_F1_357 , Final_F1_358 , Final_F1_359 , Final_F1_360 , Final_F1_361 , Final_F1_362 , Final_F1_363 , Final_F1_364 , Final_F1_365 , Final_F1_366 , Final_F1_367 , Final_F1_368 , Final_F1_369 , Final_F1_370 , Final_F1_371 , Final_F1_372 , Final_F1_373 , Final_F1_374 , Final_F1_375 , Final_F1_376 , Final_F1_377 , Final_F1_378 , Final_F1_379 , Final_F1_380 , Final_F1_381 , Final_F1_382 , Final_F1_383 , Final_F1_384 , Final_F1_385 , Final_F1_386 , Final_F1_387 , Final_F1_388 , Final_F1_389 , Final_F1_390 , Final_F1_391 , Final_F1_392 , Final_F1_393 , Final_F1_394 , Final_F1_395 , Final_F1_396 , Final_F1_397 , Final_F1_398 , Final_F1_399 , Final_F1_400 , Final_F1_401 , Final_F1_402 , Final_F1_403 , Final_F1_404 , Final_F1_405 , Final_F1_406 , Final_F1_407 , Final_F1_408 , Final_F1_409 , Final_F1_410 , Final_F1_411 , Final_F1_412 , Final_F1_413 , Final_F1_414 , Final_F1_415 , Final_F1_416 , Final_F1_417 , Final_F1_418 , Final_F1_419 , Final_F1_420 , Final_F1_421 , Final_F1_422 , Final_F1_423 , Final_F1_424 , Final_F1_425 , Final_F1_426 , Final_F1_427 , Final_F1_428 , Final_F1_429 , Final_F1_430 , Final_F1_431 , Final_F1_432 , Final_F1_433 , Final_F1_434 , Final_F1_435 , Final_F1_436 , Final_F1_437 , Final_F1_438 , Final_F1_439 , Final_F1_440 , Final_F1_441 , Final_F1_442 , Final_F1_443 , Final_F1_444 , Final_F1_445 , Final_F1_446 , Final_F1_447 , Final_F1_448 , Final_F1_449 , Final_F1_450 , Final_F1_451 , Final_F1_452 , Final_F1_453 , Final_F1_454 , Final_F1_455 , Final_F1_456 , Final_F1_457 , Final_F1_458 , Final_F1_459 , Final_F1_460 , Final_F1_461 , Final_F1_462 , Final_F1_463 , Final_F1_464 , Final_F1_465 , Final_F1_466 , Final_F1_467 , Final_F1_468 , Final_F1_469 , Final_F1_470 , Final_F1_471 , Final_F1_472 , Final_F1_473 , Final_F1_474 , Final_F1_475 , Final_F1_476 , Final_F1_477 , Final_F1_478 , Final_F1_479 , Final_F1_480 , Final_F1_481 , Final_F1_482 , Final_F1_483 , Final_F1_484 , Final_F1_485 , Final_F1_486 , Final_F1_487 , Final_F1_488 , Final_F1_489 , Final_F1_490 , Final_F1_491 , Final_F1_492 , Final_F1_493 , Final_F1_494 , Final_F1_495 , Final_F1_496 , Final_F1_497 , Final_F1_498 , Final_F1_499 , Final_F1_500 , Final_F1_501 , Final_F1_502 , Final_F1_503 , Final_F1_504 , Final_F1_505 , Final_F1_506 , Final_F1_507 , Final_F1_508 , Final_F1_509 , Final_F1_510 , Final_F1_511 , Final_F1_512 , Final_F1_513 , Final_F1_514 , Final_F1_515 , Final_F1_516 , Final_F1_517 , Final_F1_518 , Final_F1_519 , Final_F1_520 , Final_F1_521 , Final_F1_522 , Final_F1_523 , Final_F1_524 , Final_F1_525 , Final_F1_526 , Final_F1_527 , Final_F1_528 , Final_F1_529 , Final_F1_530 , Final_F1_531 , Final_F1_532 , Final_F1_533 , Final_F1_534 , Final_F1_535 , Final_F1_536 , Final_F1_537 , Final_F1_538 , Final_F1_539 , Final_F1_540 , Final_F1_541 , Final_F1_542 , Final_F1_543 , Final_F1_544 , Final_F1_545 , Final_F1_546 , Final_F1_547 , Final_F1_548 , Final_F1_549 , Final_F1_550 , Final_F1_551 , Final_F1_552 , Final_F1_553 , Final_F1_554 , Final_F1_555 , Final_F1_556 , Final_F1_557 , Final_F1_558 , Final_F1_559 , Final_F1_560 , Final_F1_561 , Final_F1_562 , Final_F1_563 , Final_F1_564 , Final_F1_565 , Final_F1_566 , Final_F1_567 , Final_F1_568 , Final_F1_569 , Final_F1_570 , Final_F1_571 , Final_F1_572 , Final_F1_573 , Final_F1_574 , Final_F1_575 ;
input wire [65:0] Final_F2_0, Final_F2_1 , Final_F2_2 , Final_F2_3 , Final_F2_4 , Final_F2_5 , Final_F2_6 , Final_F2_7 , Final_F2_8 , Final_F2_9 , Final_F2_10 , Final_F2_11 , Final_F2_12 , Final_F2_13 , Final_F2_14 , Final_F2_15 , Final_F2_16 , Final_F2_17 , Final_F2_18 , Final_F2_19 , Final_F2_20 , Final_F2_21 , Final_F2_22 , Final_F2_23 , Final_F2_24 , Final_F2_25 , Final_F2_26 , Final_F2_27 , Final_F2_28 , Final_F2_29 , Final_F2_30 , Final_F2_31 , Final_F2_32 , Final_F2_33 , Final_F2_34 , Final_F2_35 , Final_F2_36 , Final_F2_37 , Final_F2_38 , Final_F2_39 , Final_F2_40 , Final_F2_41 , Final_F2_42 , Final_F2_43 , Final_F2_44 , Final_F2_45 , Final_F2_46 , Final_F2_47 , Final_F2_48 , Final_F2_49 , Final_F2_50 , Final_F2_51 , Final_F2_52 , Final_F2_53 , Final_F2_54 , Final_F2_55 , Final_F2_56 , Final_F2_57 , Final_F2_58 , Final_F2_59 , Final_F2_60 , Final_F2_61 , Final_F2_62 , Final_F2_63 , Final_F2_64 , Final_F2_65 , Final_F2_66 , Final_F2_67 , Final_F2_68 , Final_F2_69 , Final_F2_70 , Final_F2_71 , Final_F2_72 , Final_F2_73 , Final_F2_74 , Final_F2_75 , Final_F2_76 , Final_F2_77 , Final_F2_78 , Final_F2_79 , Final_F2_80 , Final_F2_81 , Final_F2_82 , Final_F2_83 , Final_F2_84 , Final_F2_85 , Final_F2_86 , Final_F2_87 , Final_F2_88 , Final_F2_89 , Final_F2_90 , Final_F2_91 , Final_F2_92 , Final_F2_93 , Final_F2_94 , Final_F2_95 , Final_F2_96 , Final_F2_97 , Final_F2_98 , Final_F2_99 , Final_F2_100 , Final_F2_101 , Final_F2_102 , Final_F2_103 , Final_F2_104 , Final_F2_105 , Final_F2_106 , Final_F2_107 , Final_F2_108 , Final_F2_109 , Final_F2_110 , Final_F2_111 , Final_F2_112 , Final_F2_113 , Final_F2_114 , Final_F2_115 , Final_F2_116 , Final_F2_117 , Final_F2_118 , Final_F2_119 , Final_F2_120 , Final_F2_121 , Final_F2_122 , Final_F2_123 , Final_F2_124 , Final_F2_125 , Final_F2_126 , Final_F2_127 , Final_F2_128 , Final_F2_129 , Final_F2_130 , Final_F2_131 , Final_F2_132 , Final_F2_133 , Final_F2_134 , Final_F2_135 , Final_F2_136 , Final_F2_137 , Final_F2_138 , Final_F2_139 , Final_F2_140 , Final_F2_141 , Final_F2_142 , Final_F2_143 , Final_F2_144 , Final_F2_145 , Final_F2_146 , Final_F2_147 , Final_F2_148 , Final_F2_149 , Final_F2_150 , Final_F2_151 , Final_F2_152 , Final_F2_153 , Final_F2_154 , Final_F2_155 , Final_F2_156 , Final_F2_157 , Final_F2_158 , Final_F2_159 , Final_F2_160 , Final_F2_161 , Final_F2_162 , Final_F2_163 , Final_F2_164 , Final_F2_165 , Final_F2_166 , Final_F2_167 , Final_F2_168 , Final_F2_169 , Final_F2_170 , Final_F2_171 , Final_F2_172 , Final_F2_173 , Final_F2_174 , Final_F2_175 , Final_F2_176 , Final_F2_177 , Final_F2_178 , Final_F2_179 , Final_F2_180 , Final_F2_181 , Final_F2_182 , Final_F2_183 , Final_F2_184 , Final_F2_185 , Final_F2_186 , Final_F2_187 , Final_F2_188 , Final_F2_189 , Final_F2_190 , Final_F2_191 , Final_F2_192 , Final_F2_193 , Final_F2_194 , Final_F2_195 , Final_F2_196 , Final_F2_197 , Final_F2_198 , Final_F2_199 , Final_F2_200 , Final_F2_201 , Final_F2_202 , Final_F2_203 , Final_F2_204 , Final_F2_205 , Final_F2_206 , Final_F2_207 , Final_F2_208 , Final_F2_209 , Final_F2_210 , Final_F2_211 , Final_F2_212 , Final_F2_213 , Final_F2_214 , Final_F2_215 , Final_F2_216 , Final_F2_217 , Final_F2_218 , Final_F2_219 , Final_F2_220 , Final_F2_221 , Final_F2_222 , Final_F2_223 , Final_F2_224 , Final_F2_225 , Final_F2_226 , Final_F2_227 , Final_F2_228 , Final_F2_229 , Final_F2_230 , Final_F2_231 , Final_F2_232 , Final_F2_233 , Final_F2_234 , Final_F2_235 , Final_F2_236 , Final_F2_237 , Final_F2_238 , Final_F2_239 , Final_F2_240 , Final_F2_241 , Final_F2_242 , Final_F2_243 , Final_F2_244 , Final_F2_245 , Final_F2_246 , Final_F2_247 , Final_F2_248 , Final_F2_249 , Final_F2_250 , Final_F2_251 , Final_F2_252 , Final_F2_253 , Final_F2_254 , Final_F2_255 , Final_F2_256 , Final_F2_257 , Final_F2_258 , Final_F2_259 , Final_F2_260 , Final_F2_261 , Final_F2_262 , Final_F2_263 , Final_F2_264 , Final_F2_265 , Final_F2_266 , Final_F2_267 , Final_F2_268 , Final_F2_269 , Final_F2_270 , Final_F2_271 , Final_F2_272 , Final_F2_273 , Final_F2_274 , Final_F2_275 , Final_F2_276 , Final_F2_277 , Final_F2_278 , Final_F2_279 , Final_F2_280 , Final_F2_281 , Final_F2_282 , Final_F2_283 , Final_F2_284 , Final_F2_285 , Final_F2_286 , Final_F2_287 , Final_F2_288 , Final_F2_289 , Final_F2_290 , Final_F2_291 , Final_F2_292 , Final_F2_293 , Final_F2_294 , Final_F2_295 , Final_F2_296 , Final_F2_297 , Final_F2_298 , Final_F2_299 , Final_F2_300 , Final_F2_301 , Final_F2_302 , Final_F2_303 , Final_F2_304 , Final_F2_305 , Final_F2_306 , Final_F2_307 , Final_F2_308 , Final_F2_309 , Final_F2_310 , Final_F2_311 , Final_F2_312 , Final_F2_313 , Final_F2_314 , Final_F2_315 , Final_F2_316 , Final_F2_317 , Final_F2_318 , Final_F2_319 , Final_F2_320 , Final_F2_321 , Final_F2_322 , Final_F2_323 , Final_F2_324 , Final_F2_325 , Final_F2_326 , Final_F2_327 , Final_F2_328 , Final_F2_329 , Final_F2_330 , Final_F2_331 , Final_F2_332 , Final_F2_333 , Final_F2_334 , Final_F2_335 , Final_F2_336 , Final_F2_337 , Final_F2_338 , Final_F2_339 , Final_F2_340 , Final_F2_341 , Final_F2_342 , Final_F2_343 , Final_F2_344 , Final_F2_345 , Final_F2_346 , Final_F2_347 , Final_F2_348 , Final_F2_349 , Final_F2_350 , Final_F2_351 , Final_F2_352 , Final_F2_353 , Final_F2_354 , Final_F2_355 , Final_F2_356 , Final_F2_357 , Final_F2_358 , Final_F2_359 , Final_F2_360 , Final_F2_361 , Final_F2_362 , Final_F2_363 , Final_F2_364 , Final_F2_365 , Final_F2_366 , Final_F2_367 , Final_F2_368 , Final_F2_369 , Final_F2_370 , Final_F2_371 , Final_F2_372 , Final_F2_373 , Final_F2_374 , Final_F2_375 , Final_F2_376 , Final_F2_377 , Final_F2_378 , Final_F2_379 , Final_F2_380 , Final_F2_381 , Final_F2_382 , Final_F2_383 , Final_F2_384 , Final_F2_385 , Final_F2_386 , Final_F2_387 , Final_F2_388 , Final_F2_389 , Final_F2_390 , Final_F2_391 , Final_F2_392 , Final_F2_393 , Final_F2_394 , Final_F2_395 , Final_F2_396 , Final_F2_397 , Final_F2_398 , Final_F2_399 , Final_F2_400 , Final_F2_401 , Final_F2_402 , Final_F2_403 , Final_F2_404 , Final_F2_405 , Final_F2_406 , Final_F2_407 , Final_F2_408 , Final_F2_409 , Final_F2_410 , Final_F2_411 , Final_F2_412 , Final_F2_413 , Final_F2_414 , Final_F2_415 , Final_F2_416 , Final_F2_417 , Final_F2_418 , Final_F2_419 , Final_F2_420 , Final_F2_421 , Final_F2_422 , Final_F2_423 , Final_F2_424 , Final_F2_425 , Final_F2_426 , Final_F2_427 , Final_F2_428 , Final_F2_429 , Final_F2_430 , Final_F2_431 , Final_F2_432 , Final_F2_433 , Final_F2_434 , Final_F2_435 , Final_F2_436 , Final_F2_437 , Final_F2_438 , Final_F2_439 , Final_F2_440 , Final_F2_441 , Final_F2_442 , Final_F2_443 , Final_F2_444 , Final_F2_445 , Final_F2_446 , Final_F2_447 , Final_F2_448 , Final_F2_449 , Final_F2_450 , Final_F2_451 , Final_F2_452 , Final_F2_453 , Final_F2_454 , Final_F2_455 , Final_F2_456 , Final_F2_457 , Final_F2_458 , Final_F2_459 , Final_F2_460 , Final_F2_461 , Final_F2_462 , Final_F2_463 , Final_F2_464 , Final_F2_465 , Final_F2_466 , Final_F2_467 , Final_F2_468 , Final_F2_469 , Final_F2_470 , Final_F2_471 , Final_F2_472 , Final_F2_473 , Final_F2_474 , Final_F2_475 , Final_F2_476 , Final_F2_477 , Final_F2_478 , Final_F2_479 , Final_F2_480 , Final_F2_481 , Final_F2_482 , Final_F2_483 , Final_F2_484 , Final_F2_485 , Final_F2_486 , Final_F2_487 , Final_F2_488 , Final_F2_489 , Final_F2_490 , Final_F2_491 , Final_F2_492 , Final_F2_493 , Final_F2_494 , Final_F2_495 , Final_F2_496 , Final_F2_497 , Final_F2_498 , Final_F2_499 , Final_F2_500 , Final_F2_501 , Final_F2_502 , Final_F2_503 , Final_F2_504 , Final_F2_505 , Final_F2_506 , Final_F2_507 , Final_F2_508 , Final_F2_509 , Final_F2_510 , Final_F2_511 , Final_F2_512 , Final_F2_513 , Final_F2_514 , Final_F2_515 , Final_F2_516 , Final_F2_517 , Final_F2_518 , Final_F2_519 , Final_F2_520 , Final_F2_521 , Final_F2_522 , Final_F2_523 , Final_F2_524 , Final_F2_525 , Final_F2_526 , Final_F2_527 , Final_F2_528 , Final_F2_529 , Final_F2_530 , Final_F2_531 , Final_F2_532 , Final_F2_533 , Final_F2_534 , Final_F2_535 , Final_F2_536 , Final_F2_537 , Final_F2_538 , Final_F2_539 , Final_F2_540 , Final_F2_541 , Final_F2_542 , Final_F2_543 , Final_F2_544 , Final_F2_545 , Final_F2_546 , Final_F2_547 , Final_F2_548 , Final_F2_549 , Final_F2_550 , Final_F2_551 , Final_F2_552 , Final_F2_553 , Final_F2_554 , Final_F2_555 , Final_F2_556 , Final_F2_557 , Final_F2_558 , Final_F2_559 , Final_F2_560 , Final_F2_561 , Final_F2_562 , Final_F2_563 , Final_F2_564 , Final_F2_565 , Final_F2_566 , Final_F2_567 , Final_F2_568 , Final_F2_569 , Final_F2_570 , Final_F2_571 , Final_F2_572 , Final_F2_573 , Final_F2_574 , Final_F2_575 ;
input wire [65:0] Final_F3_0, Final_F3_1 , Final_F3_2 , Final_F3_3 , Final_F3_4 , Final_F3_5 , Final_F3_6 , Final_F3_7 , Final_F3_8 , Final_F3_9 , Final_F3_10 , Final_F3_11 , Final_F3_12 , Final_F3_13 , Final_F3_14 , Final_F3_15 , Final_F3_16 , Final_F3_17 , Final_F3_18 , Final_F3_19 , Final_F3_20 , Final_F3_21 , Final_F3_22 , Final_F3_23 , Final_F3_24 , Final_F3_25 , Final_F3_26 , Final_F3_27 , Final_F3_28 , Final_F3_29 , Final_F3_30 , Final_F3_31 , Final_F3_32 , Final_F3_33 , Final_F3_34 , Final_F3_35 , Final_F3_36 , Final_F3_37 , Final_F3_38 , Final_F3_39 , Final_F3_40 , Final_F3_41 , Final_F3_42 , Final_F3_43 , Final_F3_44 , Final_F3_45 , Final_F3_46 , Final_F3_47 , Final_F3_48 , Final_F3_49 , Final_F3_50 , Final_F3_51 , Final_F3_52 , Final_F3_53 , Final_F3_54 , Final_F3_55 , Final_F3_56 , Final_F3_57 , Final_F3_58 , Final_F3_59 , Final_F3_60 , Final_F3_61 , Final_F3_62 , Final_F3_63 , Final_F3_64 , Final_F3_65 , Final_F3_66 , Final_F3_67 , Final_F3_68 , Final_F3_69 , Final_F3_70 , Final_F3_71 , Final_F3_72 , Final_F3_73 , Final_F3_74 , Final_F3_75 , Final_F3_76 , Final_F3_77 , Final_F3_78 , Final_F3_79 , Final_F3_80 , Final_F3_81 , Final_F3_82 , Final_F3_83 , Final_F3_84 , Final_F3_85 , Final_F3_86 , Final_F3_87 , Final_F3_88 , Final_F3_89 , Final_F3_90 , Final_F3_91 , Final_F3_92 , Final_F3_93 , Final_F3_94 , Final_F3_95 , Final_F3_96 , Final_F3_97 , Final_F3_98 , Final_F3_99 , Final_F3_100 , Final_F3_101 , Final_F3_102 , Final_F3_103 , Final_F3_104 , Final_F3_105 , Final_F3_106 , Final_F3_107 , Final_F3_108 , Final_F3_109 , Final_F3_110 , Final_F3_111 , Final_F3_112 , Final_F3_113 , Final_F3_114 , Final_F3_115 , Final_F3_116 , Final_F3_117 , Final_F3_118 , Final_F3_119 , Final_F3_120 , Final_F3_121 , Final_F3_122 , Final_F3_123 , Final_F3_124 , Final_F3_125 , Final_F3_126 , Final_F3_127 , Final_F3_128 , Final_F3_129 , Final_F3_130 , Final_F3_131 , Final_F3_132 , Final_F3_133 , Final_F3_134 , Final_F3_135 , Final_F3_136 , Final_F3_137 , Final_F3_138 , Final_F3_139 , Final_F3_140 , Final_F3_141 , Final_F3_142 , Final_F3_143 , Final_F3_144 , Final_F3_145 , Final_F3_146 , Final_F3_147 , Final_F3_148 , Final_F3_149 , Final_F3_150 , Final_F3_151 , Final_F3_152 , Final_F3_153 , Final_F3_154 , Final_F3_155 , Final_F3_156 , Final_F3_157 , Final_F3_158 , Final_F3_159 , Final_F3_160 , Final_F3_161 , Final_F3_162 , Final_F3_163 , Final_F3_164 , Final_F3_165 , Final_F3_166 , Final_F3_167 , Final_F3_168 , Final_F3_169 , Final_F3_170 , Final_F3_171 , Final_F3_172 , Final_F3_173 , Final_F3_174 , Final_F3_175 , Final_F3_176 , Final_F3_177 , Final_F3_178 , Final_F3_179 , Final_F3_180 , Final_F3_181 , Final_F3_182 , Final_F3_183 , Final_F3_184 , Final_F3_185 , Final_F3_186 , Final_F3_187 , Final_F3_188 , Final_F3_189 , Final_F3_190 , Final_F3_191 , Final_F3_192 , Final_F3_193 , Final_F3_194 , Final_F3_195 , Final_F3_196 , Final_F3_197 , Final_F3_198 , Final_F3_199 , Final_F3_200 , Final_F3_201 , Final_F3_202 , Final_F3_203 , Final_F3_204 , Final_F3_205 , Final_F3_206 , Final_F3_207 , Final_F3_208 , Final_F3_209 , Final_F3_210 , Final_F3_211 , Final_F3_212 , Final_F3_213 , Final_F3_214 , Final_F3_215 , Final_F3_216 , Final_F3_217 , Final_F3_218 , Final_F3_219 , Final_F3_220 , Final_F3_221 , Final_F3_222 , Final_F3_223 , Final_F3_224 , Final_F3_225 , Final_F3_226 , Final_F3_227 , Final_F3_228 , Final_F3_229 , Final_F3_230 , Final_F3_231 , Final_F3_232 , Final_F3_233 , Final_F3_234 , Final_F3_235 , Final_F3_236 , Final_F3_237 , Final_F3_238 , Final_F3_239 , Final_F3_240 , Final_F3_241 , Final_F3_242 , Final_F3_243 , Final_F3_244 , Final_F3_245 , Final_F3_246 , Final_F3_247 , Final_F3_248 , Final_F3_249 , Final_F3_250 , Final_F3_251 , Final_F3_252 , Final_F3_253 , Final_F3_254 , Final_F3_255 , Final_F3_256 , Final_F3_257 , Final_F3_258 , Final_F3_259 , Final_F3_260 , Final_F3_261 , Final_F3_262 , Final_F3_263 , Final_F3_264 , Final_F3_265 , Final_F3_266 , Final_F3_267 , Final_F3_268 , Final_F3_269 , Final_F3_270 , Final_F3_271 , Final_F3_272 , Final_F3_273 , Final_F3_274 , Final_F3_275 , Final_F3_276 , Final_F3_277 , Final_F3_278 , Final_F3_279 , Final_F3_280 , Final_F3_281 , Final_F3_282 , Final_F3_283 , Final_F3_284 , Final_F3_285 , Final_F3_286 , Final_F3_287 , Final_F3_288 , Final_F3_289 , Final_F3_290 , Final_F3_291 , Final_F3_292 , Final_F3_293 , Final_F3_294 , Final_F3_295 , Final_F3_296 , Final_F3_297 , Final_F3_298 , Final_F3_299 , Final_F3_300 , Final_F3_301 , Final_F3_302 , Final_F3_303 , Final_F3_304 , Final_F3_305 , Final_F3_306 , Final_F3_307 , Final_F3_308 , Final_F3_309 , Final_F3_310 , Final_F3_311 , Final_F3_312 , Final_F3_313 , Final_F3_314 , Final_F3_315 , Final_F3_316 , Final_F3_317 , Final_F3_318 , Final_F3_319 , Final_F3_320 , Final_F3_321 , Final_F3_322 , Final_F3_323 , Final_F3_324 , Final_F3_325 , Final_F3_326 , Final_F3_327 , Final_F3_328 , Final_F3_329 , Final_F3_330 , Final_F3_331 , Final_F3_332 , Final_F3_333 , Final_F3_334 , Final_F3_335 , Final_F3_336 , Final_F3_337 , Final_F3_338 , Final_F3_339 , Final_F3_340 , Final_F3_341 , Final_F3_342 , Final_F3_343 , Final_F3_344 , Final_F3_345 , Final_F3_346 , Final_F3_347 , Final_F3_348 , Final_F3_349 , Final_F3_350 , Final_F3_351 , Final_F3_352 , Final_F3_353 , Final_F3_354 , Final_F3_355 , Final_F3_356 , Final_F3_357 , Final_F3_358 , Final_F3_359 , Final_F3_360 , Final_F3_361 , Final_F3_362 , Final_F3_363 , Final_F3_364 , Final_F3_365 , Final_F3_366 , Final_F3_367 , Final_F3_368 , Final_F3_369 , Final_F3_370 , Final_F3_371 , Final_F3_372 , Final_F3_373 , Final_F3_374 , Final_F3_375 , Final_F3_376 , Final_F3_377 , Final_F3_378 , Final_F3_379 , Final_F3_380 , Final_F3_381 , Final_F3_382 , Final_F3_383 , Final_F3_384 , Final_F3_385 , Final_F3_386 , Final_F3_387 , Final_F3_388 , Final_F3_389 , Final_F3_390 , Final_F3_391 , Final_F3_392 , Final_F3_393 , Final_F3_394 , Final_F3_395 , Final_F3_396 , Final_F3_397 , Final_F3_398 , Final_F3_399 , Final_F3_400 , Final_F3_401 , Final_F3_402 , Final_F3_403 , Final_F3_404 , Final_F3_405 , Final_F3_406 , Final_F3_407 , Final_F3_408 , Final_F3_409 , Final_F3_410 , Final_F3_411 , Final_F3_412 , Final_F3_413 , Final_F3_414 , Final_F3_415 , Final_F3_416 , Final_F3_417 , Final_F3_418 , Final_F3_419 , Final_F3_420 , Final_F3_421 , Final_F3_422 , Final_F3_423 , Final_F3_424 , Final_F3_425 , Final_F3_426 , Final_F3_427 , Final_F3_428 , Final_F3_429 , Final_F3_430 , Final_F3_431 , Final_F3_432 , Final_F3_433 , Final_F3_434 , Final_F3_435 , Final_F3_436 , Final_F3_437 , Final_F3_438 , Final_F3_439 , Final_F3_440 , Final_F3_441 , Final_F3_442 , Final_F3_443 , Final_F3_444 , Final_F3_445 , Final_F3_446 , Final_F3_447 , Final_F3_448 , Final_F3_449 , Final_F3_450 , Final_F3_451 , Final_F3_452 , Final_F3_453 , Final_F3_454 , Final_F3_455 , Final_F3_456 , Final_F3_457 , Final_F3_458 , Final_F3_459 , Final_F3_460 , Final_F3_461 , Final_F3_462 , Final_F3_463 , Final_F3_464 , Final_F3_465 , Final_F3_466 , Final_F3_467 , Final_F3_468 , Final_F3_469 , Final_F3_470 , Final_F3_471 , Final_F3_472 , Final_F3_473 , Final_F3_474 , Final_F3_475 , Final_F3_476 , Final_F3_477 , Final_F3_478 , Final_F3_479 , Final_F3_480 , Final_F3_481 , Final_F3_482 , Final_F3_483 , Final_F3_484 , Final_F3_485 , Final_F3_486 , Final_F3_487 , Final_F3_488 , Final_F3_489 , Final_F3_490 , Final_F3_491 , Final_F3_492 , Final_F3_493 , Final_F3_494 , Final_F3_495 , Final_F3_496 , Final_F3_497 , Final_F3_498 , Final_F3_499 , Final_F3_500 , Final_F3_501 , Final_F3_502 , Final_F3_503 , Final_F3_504 , Final_F3_505 , Final_F3_506 , Final_F3_507 , Final_F3_508 , Final_F3_509 , Final_F3_510 , Final_F3_511 , Final_F3_512 , Final_F3_513 , Final_F3_514 , Final_F3_515 , Final_F3_516 , Final_F3_517 , Final_F3_518 , Final_F3_519 , Final_F3_520 , Final_F3_521 , Final_F3_522 , Final_F3_523 , Final_F3_524 , Final_F3_525 , Final_F3_526 , Final_F3_527 , Final_F3_528 , Final_F3_529 , Final_F3_530 , Final_F3_531 , Final_F3_532 , Final_F3_533 , Final_F3_534 , Final_F3_535 , Final_F3_536 , Final_F3_537 , Final_F3_538 , Final_F3_539 , Final_F3_540 , Final_F3_541 , Final_F3_542 , Final_F3_543 , Final_F3_544 , Final_F3_545 , Final_F3_546 , Final_F3_547 , Final_F3_548 , Final_F3_549 , Final_F3_550 , Final_F3_551 , Final_F3_552 , Final_F3_553 , Final_F3_554 , Final_F3_555 , Final_F3_556 , Final_F3_557 , Final_F3_558 , Final_F3_559 , Final_F3_560 , Final_F3_561 , Final_F3_562 , Final_F3_563 , Final_F3_564 , Final_F3_565 , Final_F3_566 , Final_F3_567 , Final_F3_568 , Final_F3_569 , Final_F3_570 , Final_F3_571 , Final_F3_572 , Final_F3_573 , Final_F3_574 , Final_F3_575 ;
input wire [65:0] Final_F4_0, Final_F4_1 , Final_F4_2 , Final_F4_3 , Final_F4_4 , Final_F4_5 , Final_F4_6 , Final_F4_7 , Final_F4_8 , Final_F4_9 , Final_F4_10 , Final_F4_11 , Final_F4_12 , Final_F4_13 , Final_F4_14 , Final_F4_15 , Final_F4_16 , Final_F4_17 , Final_F4_18 , Final_F4_19 , Final_F4_20 , Final_F4_21 , Final_F4_22 , Final_F4_23 , Final_F4_24 , Final_F4_25 , Final_F4_26 , Final_F4_27 , Final_F4_28 , Final_F4_29 , Final_F4_30 , Final_F4_31 , Final_F4_32 , Final_F4_33 , Final_F4_34 , Final_F4_35 , Final_F4_36 , Final_F4_37 , Final_F4_38 , Final_F4_39 , Final_F4_40 , Final_F4_41 , Final_F4_42 , Final_F4_43 , Final_F4_44 , Final_F4_45 , Final_F4_46 , Final_F4_47 , Final_F4_48 , Final_F4_49 , Final_F4_50 , Final_F4_51 , Final_F4_52 , Final_F4_53 , Final_F4_54 , Final_F4_55 , Final_F4_56 , Final_F4_57 , Final_F4_58 , Final_F4_59 , Final_F4_60 , Final_F4_61 , Final_F4_62 , Final_F4_63 , Final_F4_64 , Final_F4_65 , Final_F4_66 , Final_F4_67 , Final_F4_68 , Final_F4_69 , Final_F4_70 , Final_F4_71 , Final_F4_72 , Final_F4_73 , Final_F4_74 , Final_F4_75 , Final_F4_76 , Final_F4_77 , Final_F4_78 , Final_F4_79 , Final_F4_80 , Final_F4_81 , Final_F4_82 , Final_F4_83 , Final_F4_84 , Final_F4_85 , Final_F4_86 , Final_F4_87 , Final_F4_88 , Final_F4_89 , Final_F4_90 , Final_F4_91 , Final_F4_92 , Final_F4_93 , Final_F4_94 , Final_F4_95 , Final_F4_96 , Final_F4_97 , Final_F4_98 , Final_F4_99 , Final_F4_100 , Final_F4_101 , Final_F4_102 , Final_F4_103 , Final_F4_104 , Final_F4_105 , Final_F4_106 , Final_F4_107 , Final_F4_108 , Final_F4_109 , Final_F4_110 , Final_F4_111 , Final_F4_112 , Final_F4_113 , Final_F4_114 , Final_F4_115 , Final_F4_116 , Final_F4_117 , Final_F4_118 , Final_F4_119 , Final_F4_120 , Final_F4_121 , Final_F4_122 , Final_F4_123 , Final_F4_124 , Final_F4_125 , Final_F4_126 , Final_F4_127 , Final_F4_128 , Final_F4_129 , Final_F4_130 , Final_F4_131 , Final_F4_132 , Final_F4_133 , Final_F4_134 , Final_F4_135 , Final_F4_136 , Final_F4_137 , Final_F4_138 , Final_F4_139 , Final_F4_140 , Final_F4_141 , Final_F4_142 , Final_F4_143 , Final_F4_144 , Final_F4_145 , Final_F4_146 , Final_F4_147 , Final_F4_148 , Final_F4_149 , Final_F4_150 , Final_F4_151 , Final_F4_152 , Final_F4_153 , Final_F4_154 , Final_F4_155 , Final_F4_156 , Final_F4_157 , Final_F4_158 , Final_F4_159 , Final_F4_160 , Final_F4_161 , Final_F4_162 , Final_F4_163 , Final_F4_164 , Final_F4_165 , Final_F4_166 , Final_F4_167 , Final_F4_168 , Final_F4_169 , Final_F4_170 , Final_F4_171 , Final_F4_172 , Final_F4_173 , Final_F4_174 , Final_F4_175 , Final_F4_176 , Final_F4_177 , Final_F4_178 , Final_F4_179 , Final_F4_180 , Final_F4_181 , Final_F4_182 , Final_F4_183 , Final_F4_184 , Final_F4_185 , Final_F4_186 , Final_F4_187 , Final_F4_188 , Final_F4_189 , Final_F4_190 , Final_F4_191 , Final_F4_192 , Final_F4_193 , Final_F4_194 , Final_F4_195 , Final_F4_196 , Final_F4_197 , Final_F4_198 , Final_F4_199 , Final_F4_200 , Final_F4_201 , Final_F4_202 , Final_F4_203 , Final_F4_204 , Final_F4_205 , Final_F4_206 , Final_F4_207 , Final_F4_208 , Final_F4_209 , Final_F4_210 , Final_F4_211 , Final_F4_212 , Final_F4_213 , Final_F4_214 , Final_F4_215 , Final_F4_216 , Final_F4_217 , Final_F4_218 , Final_F4_219 , Final_F4_220 , Final_F4_221 , Final_F4_222 , Final_F4_223 , Final_F4_224 , Final_F4_225 , Final_F4_226 , Final_F4_227 , Final_F4_228 , Final_F4_229 , Final_F4_230 , Final_F4_231 , Final_F4_232 , Final_F4_233 , Final_F4_234 , Final_F4_235 , Final_F4_236 , Final_F4_237 , Final_F4_238 , Final_F4_239 , Final_F4_240 , Final_F4_241 , Final_F4_242 , Final_F4_243 , Final_F4_244 , Final_F4_245 , Final_F4_246 , Final_F4_247 , Final_F4_248 , Final_F4_249 , Final_F4_250 , Final_F4_251 , Final_F4_252 , Final_F4_253 , Final_F4_254 , Final_F4_255 , Final_F4_256 , Final_F4_257 , Final_F4_258 , Final_F4_259 , Final_F4_260 , Final_F4_261 , Final_F4_262 , Final_F4_263 , Final_F4_264 , Final_F4_265 , Final_F4_266 , Final_F4_267 , Final_F4_268 , Final_F4_269 , Final_F4_270 , Final_F4_271 , Final_F4_272 , Final_F4_273 , Final_F4_274 , Final_F4_275 , Final_F4_276 , Final_F4_277 , Final_F4_278 , Final_F4_279 , Final_F4_280 , Final_F4_281 , Final_F4_282 , Final_F4_283 , Final_F4_284 , Final_F4_285 , Final_F4_286 , Final_F4_287 , Final_F4_288 , Final_F4_289 , Final_F4_290 , Final_F4_291 , Final_F4_292 , Final_F4_293 , Final_F4_294 , Final_F4_295 , Final_F4_296 , Final_F4_297 , Final_F4_298 , Final_F4_299 , Final_F4_300 , Final_F4_301 , Final_F4_302 , Final_F4_303 , Final_F4_304 , Final_F4_305 , Final_F4_306 , Final_F4_307 , Final_F4_308 , Final_F4_309 , Final_F4_310 , Final_F4_311 , Final_F4_312 , Final_F4_313 , Final_F4_314 , Final_F4_315 , Final_F4_316 , Final_F4_317 , Final_F4_318 , Final_F4_319 , Final_F4_320 , Final_F4_321 , Final_F4_322 , Final_F4_323 , Final_F4_324 , Final_F4_325 , Final_F4_326 , Final_F4_327 , Final_F4_328 , Final_F4_329 , Final_F4_330 , Final_F4_331 , Final_F4_332 , Final_F4_333 , Final_F4_334 , Final_F4_335 , Final_F4_336 , Final_F4_337 , Final_F4_338 , Final_F4_339 , Final_F4_340 , Final_F4_341 , Final_F4_342 , Final_F4_343 , Final_F4_344 , Final_F4_345 , Final_F4_346 , Final_F4_347 , Final_F4_348 , Final_F4_349 , Final_F4_350 , Final_F4_351 , Final_F4_352 , Final_F4_353 , Final_F4_354 , Final_F4_355 , Final_F4_356 , Final_F4_357 , Final_F4_358 , Final_F4_359 , Final_F4_360 , Final_F4_361 , Final_F4_362 , Final_F4_363 , Final_F4_364 , Final_F4_365 , Final_F4_366 , Final_F4_367 , Final_F4_368 , Final_F4_369 , Final_F4_370 , Final_F4_371 , Final_F4_372 , Final_F4_373 , Final_F4_374 , Final_F4_375 , Final_F4_376 , Final_F4_377 , Final_F4_378 , Final_F4_379 , Final_F4_380 , Final_F4_381 , Final_F4_382 , Final_F4_383 , Final_F4_384 , Final_F4_385 , Final_F4_386 , Final_F4_387 , Final_F4_388 , Final_F4_389 , Final_F4_390 , Final_F4_391 , Final_F4_392 , Final_F4_393 , Final_F4_394 , Final_F4_395 , Final_F4_396 , Final_F4_397 , Final_F4_398 , Final_F4_399 , Final_F4_400 , Final_F4_401 , Final_F4_402 , Final_F4_403 , Final_F4_404 , Final_F4_405 , Final_F4_406 , Final_F4_407 , Final_F4_408 , Final_F4_409 , Final_F4_410 , Final_F4_411 , Final_F4_412 , Final_F4_413 , Final_F4_414 , Final_F4_415 , Final_F4_416 , Final_F4_417 , Final_F4_418 , Final_F4_419 , Final_F4_420 , Final_F4_421 , Final_F4_422 , Final_F4_423 , Final_F4_424 , Final_F4_425 , Final_F4_426 , Final_F4_427 , Final_F4_428 , Final_F4_429 , Final_F4_430 , Final_F4_431 , Final_F4_432 , Final_F4_433 , Final_F4_434 , Final_F4_435 , Final_F4_436 , Final_F4_437 , Final_F4_438 , Final_F4_439 , Final_F4_440 , Final_F4_441 , Final_F4_442 , Final_F4_443 , Final_F4_444 , Final_F4_445 , Final_F4_446 , Final_F4_447 , Final_F4_448 , Final_F4_449 , Final_F4_450 , Final_F4_451 , Final_F4_452 , Final_F4_453 , Final_F4_454 , Final_F4_455 , Final_F4_456 , Final_F4_457 , Final_F4_458 , Final_F4_459 , Final_F4_460 , Final_F4_461 , Final_F4_462 , Final_F4_463 , Final_F4_464 , Final_F4_465 , Final_F4_466 , Final_F4_467 , Final_F4_468 , Final_F4_469 , Final_F4_470 , Final_F4_471 , Final_F4_472 , Final_F4_473 , Final_F4_474 , Final_F4_475 , Final_F4_476 , Final_F4_477 , Final_F4_478 , Final_F4_479 , Final_F4_480 , Final_F4_481 , Final_F4_482 , Final_F4_483 , Final_F4_484 , Final_F4_485 , Final_F4_486 , Final_F4_487 , Final_F4_488 , Final_F4_489 , Final_F4_490 , Final_F4_491 , Final_F4_492 , Final_F4_493 , Final_F4_494 , Final_F4_495 , Final_F4_496 , Final_F4_497 , Final_F4_498 , Final_F4_499 , Final_F4_500 , Final_F4_501 , Final_F4_502 , Final_F4_503 , Final_F4_504 , Final_F4_505 , Final_F4_506 , Final_F4_507 , Final_F4_508 , Final_F4_509 , Final_F4_510 , Final_F4_511 , Final_F4_512 , Final_F4_513 , Final_F4_514 , Final_F4_515 , Final_F4_516 , Final_F4_517 , Final_F4_518 , Final_F4_519 , Final_F4_520 , Final_F4_521 , Final_F4_522 , Final_F4_523 , Final_F4_524 , Final_F4_525 , Final_F4_526 , Final_F4_527 , Final_F4_528 , Final_F4_529 , Final_F4_530 , Final_F4_531 , Final_F4_532 , Final_F4_533 , Final_F4_534 , Final_F4_535 , Final_F4_536 , Final_F4_537 , Final_F4_538 , Final_F4_539 , Final_F4_540 , Final_F4_541 , Final_F4_542 , Final_F4_543 , Final_F4_544 , Final_F4_545 , Final_F4_546 , Final_F4_547 , Final_F4_548 , Final_F4_549 , Final_F4_550 , Final_F4_551 , Final_F4_552 , Final_F4_553 , Final_F4_554 , Final_F4_555 , Final_F4_556 , Final_F4_557 , Final_F4_558 , Final_F4_559 , Final_F4_560 , Final_F4_561 , Final_F4_562 , Final_F4_563 , Final_F4_564 , Final_F4_565 , Final_F4_566 , Final_F4_567 , Final_F4_568 , Final_F4_569 , Final_F4_570 , Final_F4_571 , Final_F4_572 , Final_F4_573 , Final_F4_574 , Final_F4_575 ;
 */
/* 
output wire [65:0]  REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143; 
output wire [65:0]  REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143; 
output wire [65:0]  REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143; 
output wire [65:0]  REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143; 
  */

 
//reg MAXwrite2_1 , MAXwrite2_2 , MAXwrite2_3 , MAXwrite2_4 , MAXwrite2_5 , MAXwrite2_6 , MAXwrite2_7 , MAXwrite2_8 , MAXwrite2_9 , MAXwrite2_10 , MAXwrite2_11 , MAXwrite2_12 , MAXwrite2_13 , MAXwrite2_14 , MAXwrite2_15 , MAXwrite2_16 , MAXwrite2_17 , MAXwrite2_18 , MAXwrite2_19 , MAXwrite2_20 , MAXwrite2_21 , MAXwrite2_22 , MAXwrite2_23 , MAXwrite2_24 , MAXwrite2_25 , MAXwrite2_26 , MAXwrite2_27 , MAXwrite2_28 , MAXwrite2_29 , MAXwrite2_30 , MAXwrite2_31 , MAXwrite2_32 , MAXwrite2_33 , MAXwrite2_34 , MAXwrite2_35 , MAXwrite2_36 , MAXwrite2_37 , MAXwrite2_38 , MAXwrite2_39 , MAXwrite2_40 , MAXwrite2_41 , MAXwrite2_42 , MAXwrite2_43 , MAXwrite2_44 , MAXwrite2_45 , MAXwrite2_46 , MAXwrite2_47 , MAXwrite2_48 , MAXwrite2_49 , MAXwrite2_50 , MAXwrite2_51 , MAXwrite2_52 , MAXwrite2_53 , MAXwrite2_54 , MAXwrite2_55 , MAXwrite2_56 , MAXwrite2_57 , MAXwrite2_58 , MAXwrite2_59 , MAXwrite2_60 , MAXwrite2_61 , MAXwrite2_62 , MAXwrite2_63 , MAXwrite2_64 , MAXwrite2_65 , MAXwrite2_66 , MAXwrite2_67 , MAXwrite2_68 , MAXwrite2_69 , MAXwrite2_70 , MAXwrite2_71 , MAXwrite2_72 , MAXwrite2_73 , MAXwrite2_74 , MAXwrite2_75 , MAXwrite2_76 , MAXwrite2_77 , MAXwrite2_78 , MAXwrite2_79 , MAXwrite2_80 , MAXwrite2_81 , MAXwrite2_82 , MAXwrite2_83 , MAXwrite2_84 , MAXwrite2_85 , MAXwrite2_86 , MAXwrite2_87 , MAXwrite2_88 , MAXwrite2_89 , MAXwrite2_90 , MAXwrite2_91 , MAXwrite2_92 , MAXwrite2_93 , MAXwrite2_94 , MAXwrite2_95 , MAXwrite2_96 , MAXwrite2_97 , MAXwrite2_98 , MAXwrite2_99 , MAXwrite2_100 , MAXwrite2_101 , MAXwrite2_102 , MAXwrite2_103 , MAXwrite2_104 , MAXwrite2_105 , MAXwrite2_106 , MAXwrite2_107 , MAXwrite2_108 , MAXwrite2_109 , MAXwrite2_110 , MAXwrite2_111 , MAXwrite2_112 , MAXwrite2_113 , MAXwrite2_114 , MAXwrite2_115 , MAXwrite2_116 , MAXwrite2_117 , MAXwrite2_118 , MAXwrite2_119 , MAXwrite2_120 , MAXwrite2_121 , MAXwrite2_122 , MAXwrite2_123 , MAXwrite2_124 , MAXwrite2_125 , MAXwrite2_126 , MAXwrite2_127 , MAXwrite2_128 , MAXwrite2_129 , MAXwrite2_130 , MAXwrite2_131 , MAXwrite2_132 , MAXwrite2_133 , MAXwrite2_134 , MAXwrite2_135 , MAXwrite2_136 , MAXwrite2_137 , MAXwrite2_138 , MAXwrite2_139 , MAXwrite2_140 , MAXwrite2_141 , MAXwrite2_142 , MAXwrite2_143 , MAXwrite2_144 ;



/* always @ (posedge clk)
begin
if (superADDRESS ==   2) begin  
MAXwrite2_1  <= 1; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
end

else if (superADDRESS ==   5) begin
MAXwrite2_1  <= 0; MAXwrite2_2   <= 1; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
          end 
else if (superADDRESS ==   8) begin 
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 1;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
         end 
else if (superADDRESS ==   11) begin 
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 1;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
         end 
else if (superADDRESS ==   14) begin  
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 1;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
        end 
else if (superADDRESS ==   17) begin  
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 1; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
        end 
else if (superADDRESS ==   20) begin
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 1;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
          end 
else if (superADDRESS ==   23) begin 
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 1; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
         end 
else if (superADDRESS ==   26) begin 
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 1;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
         end 
else if (superADDRESS ==   29) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 1; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
       end 
else if (superADDRESS ==   32) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 1;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
       end 
else if (superADDRESS ==   35) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 1;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
      end 
else if (superADDRESS ==   38) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 1;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
      end 
else if (superADDRESS ==   41) begin  
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 1; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
        end 
else if (superADDRESS ==   44) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 1;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
      end 
else if (superADDRESS ==   47) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 1; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
      end 
else if (superADDRESS ==   50) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 1;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
       end 
else if (superADDRESS ==   53) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 1; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
       end 
else if (superADDRESS ==   56) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 1;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
       end 
else if (superADDRESS ==   59) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 1;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
       end 
else if (superADDRESS ==   62) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 1;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
    end 
else if (superADDRESS ==   65) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 1; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
      end 
else if (superADDRESS ==   68) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 1;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
      end 
else if (superADDRESS ==   71) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 1; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
      end 
else if (superADDRESS ==   74) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 1;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
      end 
else if (superADDRESS ==   77) begin  

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 1; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;       end 
else if (superADDRESS ==   80) begin  
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 1;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;       end 
else if (superADDRESS ==   83) begin  

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 1;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;       end 
else if (superADDRESS ==   86) begin  

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 1;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;       end 
else if (superADDRESS ==   89) begin 

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 1; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;        end 
else if (superADDRESS ==   92) begin   

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 1;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   95) begin 

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 1; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;        end 
else if (superADDRESS ==   98) begin 

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 1;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;        end 
else if (superADDRESS ==   101) begin   

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 1; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   104) begin   

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 1;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   107) begin  
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 1;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;       end 
else if (superADDRESS ==   110) begin   

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 1;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   113) begin  

MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 1; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;       end 
else if (superADDRESS ==   116) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 1;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   119) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 1; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   122) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 1;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   125) begin  
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 1; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;       end 
else if (superADDRESS ==   128) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 1;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   131) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 1;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   134) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 1;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   137) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 1; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   140) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 1;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   143) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 1; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   146) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 1;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   149) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 1; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   152) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 1;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   155) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 1;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   158) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 1;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   161) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 1; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   164) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 1;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   167) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 1; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   170) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 1;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   173) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 1; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   176) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 1;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   179) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 1;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   182) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 1;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   185) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 1; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   188) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 1;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   191) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 1; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   194) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 1;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   197) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 1; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   200) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 1;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   203) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 1;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   206) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 1;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   209) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 1; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   212) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 1;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   215) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 1; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   218) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 1;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   221) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 1; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   224) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 1;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   227) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 1;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   230) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 1;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   233) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 1; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   236) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 1;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   239) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 1; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   242) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 1;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   245) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 1; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   248) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 1;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   251) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 1;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   254) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 1;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   257) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 1; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   260) begin       
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 1;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;  end 
else if (superADDRESS ==   263) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 1; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   266) begin        
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 1;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; end 
else if (superADDRESS ==   269) begin       
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 1; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;  end 
else if (superADDRESS ==   272) begin       
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 1;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;  end 
else if (superADDRESS ==   275) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 1;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   278) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 1;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   281) begin       
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 1; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;  end 
else if (superADDRESS ==   284) begin       
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 1;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;  end 
else if (superADDRESS ==   287) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 1; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   290) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 1;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   293) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 1; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   296) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 1;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   299) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 1;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   302) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 1;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   305) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 1; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   308) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 1;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   311) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 1; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   314) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 1;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   317) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 1; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   320) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 1;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   323) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 1;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   326) begin       
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 1;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;  end 
else if (superADDRESS ==   329) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 1; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   332) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 1;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   335) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 1; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   338) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 1;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   341) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 1; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   344) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 1;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   347) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 1;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   350) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 1;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   353) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 1; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   356) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 1;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   359) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 1; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   362) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 1;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   365) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 1; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   368) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 1;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   371) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 1;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   374) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 1;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   377) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 1; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   380) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 1;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   383) begin       
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 1; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;  end 
else if (superADDRESS ==   386) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 1;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   389) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 1; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   392) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 1;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   395) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 1;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   398) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 1;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   401) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 1; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   404) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 1;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   407) begin    
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 1; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;     end 
else if (superADDRESS ==   410) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 1;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;      end 
else if (superADDRESS ==   413) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 1; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   416) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 1;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   419) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 1;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   422) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 1;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   425) begin     
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 1; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0;    end 
else if (superADDRESS ==   428) begin      
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 1;  MAXwrite2_144   <= 0;   end 
else if (superADDRESS ==   431) begin   
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 1;      end 


else begin  
MAXwrite2_1  <= 0; MAXwrite2_2   <= 0; MAXwrite2_3   <= 0;  MAXwrite2_4   <= 0;  MAXwrite2_5   <= 0;  MAXwrite2_6   <= 0; MAXwrite2_7   <= 0;  MAXwrite2_8   <= 0; 
MAXwrite2_9  <= 0;  MAXwrite2_10   <= 0; MAXwrite2_11   <= 0;  MAXwrite2_12   <= 0;  MAXwrite2_13   <= 0;  MAXwrite2_14   <= 0; MAXwrite2_15   <= 0;  MAXwrite2_16   <= 0; 
MAXwrite2_17  <= 0;  MAXwrite2_18   <= 0; MAXwrite2_19   <= 0;  MAXwrite2_20   <= 0;  MAXwrite2_21   <= 0;  MAXwrite2_22   <= 0; MAXwrite2_23   <= 0;  MAXwrite2_24   <= 0; 
MAXwrite2_25  <= 0;  MAXwrite2_26   <= 0; MAXwrite2_27   <= 0;  MAXwrite2_28   <= 0;  MAXwrite2_29   <= 0;  MAXwrite2_30   <= 0; MAXwrite2_31   <= 0;  MAXwrite2_32   <= 0; 
MAXwrite2_33  <= 0;  MAXwrite2_34   <= 0; MAXwrite2_35   <= 0;  MAXwrite2_36   <= 0;  MAXwrite2_37   <= 0;  MAXwrite2_38   <= 0; MAXwrite2_39   <= 0;  MAXwrite2_40   <= 0; 
MAXwrite2_41  <= 0;  MAXwrite2_42   <= 0; MAXwrite2_43   <= 0;  MAXwrite2_44   <= 0;  MAXwrite2_45   <= 0;  MAXwrite2_46   <= 0; MAXwrite2_47   <= 0;  MAXwrite2_48   <= 0; 
MAXwrite2_49  <= 0;  MAXwrite2_50   <= 0; MAXwrite2_51   <= 0;  MAXwrite2_52   <= 0;  MAXwrite2_53   <= 0;  MAXwrite2_54   <= 0; MAXwrite2_55   <= 0;  MAXwrite2_56   <= 0; 
MAXwrite2_57  <= 0;  MAXwrite2_58   <= 0; MAXwrite2_59   <= 0;  MAXwrite2_60   <= 0;  MAXwrite2_61   <= 0;  MAXwrite2_62   <= 0; MAXwrite2_63   <= 0;  MAXwrite2_64   <= 0; 
MAXwrite2_65  <= 0;  MAXwrite2_66   <= 0; MAXwrite2_67   <= 0;  MAXwrite2_68   <= 0;  MAXwrite2_69   <= 0;  MAXwrite2_70   <= 0; MAXwrite2_71   <= 0;  MAXwrite2_72   <= 0; 
MAXwrite2_73  <= 0;  MAXwrite2_74   <= 0; MAXwrite2_75   <= 0;  MAXwrite2_76   <= 0;  MAXwrite2_77   <= 0;  MAXwrite2_78   <= 0; MAXwrite2_79   <= 0;  MAXwrite2_80   <= 0; 
MAXwrite2_81  <= 0;  MAXwrite2_82   <= 0; MAXwrite2_83   <= 0;  MAXwrite2_84   <= 0;  MAXwrite2_85   <= 0;  MAXwrite2_86   <= 0; MAXwrite2_87   <= 0;  MAXwrite2_88   <= 0; 
MAXwrite2_89  <= 0;  MAXwrite2_90   <= 0; MAXwrite2_91   <= 0;  MAXwrite2_92   <= 0;  MAXwrite2_93   <= 0;  MAXwrite2_94   <= 0; MAXwrite2_95   <= 0;  MAXwrite2_96   <= 0; 
MAXwrite2_97  <= 0;  MAXwrite2_98   <= 0; MAXwrite2_99   <= 0;  MAXwrite2_100   <= 0;  MAXwrite2_101   <= 0;  MAXwrite2_102   <= 0; MAXwrite2_103   <= 0;  MAXwrite2_104   <= 0; 
MAXwrite2_105  <= 0;  MAXwrite2_106   <= 0; MAXwrite2_107   <= 0;  MAXwrite2_108   <= 0;  MAXwrite2_109   <= 0;  MAXwrite2_110   <= 0; MAXwrite2_111   <= 0;  MAXwrite2_112   <= 0; 
MAXwrite2_113  <= 0;  MAXwrite2_114   <= 0; MAXwrite2_115   <= 0;  MAXwrite2_116   <= 0;  MAXwrite2_117   <= 0;  MAXwrite2_118   <= 0; MAXwrite2_119   <= 0;  MAXwrite2_120   <= 0; 
MAXwrite2_121  <= 0;  MAXwrite2_122   <= 0; MAXwrite2_123   <= 0;  MAXwrite2_124   <= 0;  MAXwrite2_125   <= 0;  MAXwrite2_126   <= 0; MAXwrite2_127   <= 0;  MAXwrite2_128   <= 0; 
MAXwrite2_129  <= 0;  MAXwrite2_130   <= 0; MAXwrite2_131   <= 0;  MAXwrite2_132   <= 0;  MAXwrite2_133   <= 0;  MAXwrite2_134   <= 0; MAXwrite2_135   <= 0;  MAXwrite2_136   <= 0; 
MAXwrite2_137  <= 0;  MAXwrite2_138   <= 0; MAXwrite2_139   <= 0;  MAXwrite2_140   <= 0;  MAXwrite2_141   <= 0;  MAXwrite2_142   <= 0; MAXwrite2_143   <= 0;  MAXwrite2_144   <= 0; 
 end

end

 */



wire [65:0]  /* SuperMuxOut_F1_1, SuperMuxOut_F1_2, SuperMuxOut_F1_3, SuperMuxOut_F1_4 , */ CompOut_F1;
wire [65:0] /*  SuperMuxOut_F2_1, SuperMuxOut_F2_2, SuperMuxOut_F2_3, SuperMuxOut_F2_4 ,  */ CompOut_F2;
wire [65:0] /*  SuperMuxOut_F3_1, SuperMuxOut_F3_2, SuperMuxOut_F3_3, SuperMuxOut_F3_4 ,  */ CompOut_F3;
wire [65:0]  /* SuperMuxOut_F4_1, SuperMuxOut_F4_2, SuperMuxOut_F4_3, SuperMuxOut_F4_4 ,  */ CompOut_F4;


//COUNTER_LAYER_433_cycles MAX1TheCounter(clk,superADDRESS, MAX1LayerStart,MAX1LayerFinish );


//1//

/*
SUPERMUXMODULE_MAXPOOL1_2by2_340 F1_1_1_1 
( Final_F1_0 , Final_F1_2 , Final_F1_4 , Final_F1_6 , Final_F1_8 , Final_F1_10 , Final_F1_12 , Final_F1_14 , Final_F1_16 , Final_F1_18 , Final_F1_20 , Final_F1_22
, Final_F1_48 , Final_F1_50 , Final_F1_52 , Final_F1_54 , Final_F1_56 , Final_F1_58 , Final_F1_60 , Final_F1_62 , Final_F1_64 , Final_F1_66 , Final_F1_68 , Final_F1_70
, Final_F1_96 , Final_F1_98 , Final_F1_100 , Final_F1_102 , Final_F1_104 , Final_F1_106 , Final_F1_108 , Final_F1_110 , Final_F1_112 , Final_F1_114 , Final_F1_116 , Final_F1_118
, Final_F1_144 , Final_F1_146 , Final_F1_148 , Final_F1_150 , Final_F1_152 , Final_F1_154 , Final_F1_156 , Final_F1_158 , Final_F1_160 , Final_F1_162 , Final_F1_164 , Final_F1_166
, Final_F1_192 , Final_F1_194 , Final_F1_196 , Final_F1_198 , Final_F1_200 , Final_F1_202 , Final_F1_204 , Final_F1_206 , Final_F1_208 , Final_F1_210 , Final_F1_212 , Final_F1_214
, Final_F1_240 , Final_F1_242 , Final_F1_244 , Final_F1_246 , Final_F1_248 , Final_F1_250 , Final_F1_252 , Final_F1_254 , Final_F1_256 , Final_F1_258 , Final_F1_260 , Final_F1_262
, Final_F1_288 , Final_F1_290 , Final_F1_292 , Final_F1_294 , Final_F1_296 , Final_F1_298 , Final_F1_300 , Final_F1_302 , Final_F1_304 , Final_F1_306 , Final_F1_308 , Final_F1_310
, Final_F1_336 , Final_F1_338 , Final_F1_340 , Final_F1_342 , Final_F1_344 , Final_F1_346 , Final_F1_348 , Final_F1_350 , Final_F1_352 , Final_F1_354 , Final_F1_356 , Final_F1_358
, Final_F1_384 , Final_F1_386 , Final_F1_388 , Final_F1_390 , Final_F1_392 , Final_F1_394 , Final_F1_396 , Final_F1_398 , Final_F1_400 , Final_F1_402 , Final_F1_404 , Final_F1_406
, Final_F1_432 , Final_F1_434 , Final_F1_436 , Final_F1_438 , Final_F1_440 , Final_F1_442 , Final_F1_444 , Final_F1_446 , Final_F1_448 , Final_F1_450 , Final_F1_452 , Final_F1_454
, Final_F1_480 , Final_F1_482 , Final_F1_484 , Final_F1_486 , Final_F1_488 , Final_F1_490 , Final_F1_492 , Final_F1_494 , Final_F1_496 , Final_F1_498 , Final_F1_500 , Final_F1_502
, Final_F1_528 , Final_F1_530 , Final_F1_532 , Final_F1_534 , Final_F1_536 , Final_F1_538 , Final_F1_540 , Final_F1_542 , Final_F1_544 , Final_F1_546 , Final_F1_548 , Final_F1_550
, superADDRESS, SuperMuxOut_F1_1);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F1_1_1_2 
( Final_F1_1 , Final_F1_3 , Final_F1_5 , Final_F1_7 , Final_F1_9 , Final_F1_11 , Final_F1_13 , Final_F1_15 , Final_F1_17 , Final_F1_19 , Final_F1_21 , Final_F1_23
, Final_F1_49 , Final_F1_51 , Final_F1_53 , Final_F1_55 , Final_F1_57 , Final_F1_59 , Final_F1_61 , Final_F1_63 , Final_F1_65 , Final_F1_67 , Final_F1_69 , Final_F1_71
, Final_F1_97 , Final_F1_99 , Final_F1_101 , Final_F1_103 , Final_F1_105 , Final_F1_107 , Final_F1_109 , Final_F1_111 , Final_F1_113 , Final_F1_115 , Final_F1_117 , Final_F1_119
, Final_F1_145 , Final_F1_147 , Final_F1_149 , Final_F1_151 , Final_F1_153 , Final_F1_155 , Final_F1_157 , Final_F1_159 , Final_F1_161 , Final_F1_163 , Final_F1_165 , Final_F1_167
, Final_F1_193 , Final_F1_195 , Final_F1_197 , Final_F1_199 , Final_F1_201 , Final_F1_203 , Final_F1_205 , Final_F1_207 , Final_F1_209 , Final_F1_211 , Final_F1_213 , Final_F1_215
, Final_F1_241 , Final_F1_243 , Final_F1_245 , Final_F1_247 , Final_F1_249 , Final_F1_251 , Final_F1_253 , Final_F1_255 , Final_F1_257 , Final_F1_259 , Final_F1_261 , Final_F1_263
, Final_F1_289 , Final_F1_291 , Final_F1_293 , Final_F1_295 , Final_F1_297 , Final_F1_299 , Final_F1_301 , Final_F1_303 , Final_F1_305 , Final_F1_307 , Final_F1_309 , Final_F1_311
, Final_F1_337 , Final_F1_339 , Final_F1_341 , Final_F1_343 , Final_F1_345 , Final_F1_347 , Final_F1_349 , Final_F1_351 , Final_F1_353 , Final_F1_355 , Final_F1_357 , Final_F1_359
, Final_F1_385 , Final_F1_387 , Final_F1_389 , Final_F1_391 , Final_F1_393 , Final_F1_395 , Final_F1_397 , Final_F1_399 , Final_F1_401 , Final_F1_403 , Final_F1_405 , Final_F1_407
, Final_F1_433 , Final_F1_435 , Final_F1_437 , Final_F1_439 , Final_F1_441 , Final_F1_443 , Final_F1_445 , Final_F1_447 , Final_F1_449 , Final_F1_451 , Final_F1_453 , Final_F1_455
, Final_F1_481 , Final_F1_483 , Final_F1_485 , Final_F1_487 , Final_F1_489 , Final_F1_491 , Final_F1_493 , Final_F1_495 , Final_F1_497 , Final_F1_499 , Final_F1_501 , Final_F1_503
, Final_F1_529 , Final_F1_531 , Final_F1_533 , Final_F1_535 , Final_F1_537 , Final_F1_539 , Final_F1_541 , Final_F1_543 , Final_F1_545 , Final_F1_547 , Final_F1_549 , Final_F1_551
, superADDRESS, SuperMuxOut_F1_2);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F1_1_1_3 
( Final_F1_24 , Final_F1_26 , Final_F1_28 , Final_F1_30 , Final_F1_32 , Final_F1_34 , Final_F1_36 , Final_F1_38 , Final_F1_40 , Final_F1_42 , Final_F1_44 , Final_F1_46
, Final_F1_72 , Final_F1_74 , Final_F1_76 , Final_F1_78 , Final_F1_80 , Final_F1_82 , Final_F1_84 , Final_F1_86 , Final_F1_88 , Final_F1_90 , Final_F1_92 , Final_F1_94
, Final_F1_120 , Final_F1_122 , Final_F1_124 , Final_F1_126 , Final_F1_128 , Final_F1_130 , Final_F1_132 , Final_F1_134 , Final_F1_136 , Final_F1_138 , Final_F1_140 , Final_F1_142
, Final_F1_168 , Final_F1_170 , Final_F1_172 , Final_F1_174 , Final_F1_176 , Final_F1_178 , Final_F1_180 , Final_F1_182 , Final_F1_184 , Final_F1_186 , Final_F1_188 , Final_F1_190
, Final_F1_216 , Final_F1_218 , Final_F1_220 , Final_F1_222 , Final_F1_224 , Final_F1_226 , Final_F1_228 , Final_F1_230 , Final_F1_232 , Final_F1_234 , Final_F1_236 , Final_F1_238
, Final_F1_264 , Final_F1_266 , Final_F1_268 , Final_F1_270 , Final_F1_272 , Final_F1_274 , Final_F1_276 , Final_F1_278 , Final_F1_280 , Final_F1_282 , Final_F1_284 , Final_F1_286
, Final_F1_312 , Final_F1_314 , Final_F1_316 , Final_F1_318 , Final_F1_320 , Final_F1_322 , Final_F1_324 , Final_F1_326 , Final_F1_328 , Final_F1_330 , Final_F1_332 , Final_F1_334
, Final_F1_360 , Final_F1_362 , Final_F1_364 , Final_F1_366 , Final_F1_368 , Final_F1_370 , Final_F1_372 , Final_F1_374 , Final_F1_376 , Final_F1_378 , Final_F1_380 , Final_F1_382
, Final_F1_408 , Final_F1_410 , Final_F1_412 , Final_F1_414 , Final_F1_416 , Final_F1_418 , Final_F1_420 , Final_F1_422 , Final_F1_424 , Final_F1_426 , Final_F1_428 , Final_F1_430
, Final_F1_456 , Final_F1_458 , Final_F1_460 , Final_F1_462 , Final_F1_464 , Final_F1_466 , Final_F1_468 , Final_F1_470 , Final_F1_472 , Final_F1_474 , Final_F1_476 , Final_F1_478
, Final_F1_504 , Final_F1_506 , Final_F1_508 , Final_F1_510 , Final_F1_512 , Final_F1_514 , Final_F1_516 , Final_F1_518 , Final_F1_520 , Final_F1_522 , Final_F1_524 , Final_F1_526
, Final_F1_552 , Final_F1_554 , Final_F1_556 , Final_F1_558 , Final_F1_560 , Final_F1_562 , Final_F1_564 , Final_F1_566 , Final_F1_568 , Final_F1_570 , Final_F1_572 , Final_F1_574
, superADDRESS, SuperMuxOut_F1_3);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F1_1_1_4
( Final_F1_25 , Final_F1_27 , Final_F1_29 , Final_F1_31 , Final_F1_33 , Final_F1_35 , Final_F1_37 , Final_F1_39 , Final_F1_41 , Final_F1_43 , Final_F1_45 , Final_F1_47
, Final_F1_73 , Final_F1_75 , Final_F1_77 , Final_F1_79 , Final_F1_81 , Final_F1_83 , Final_F1_85 , Final_F1_87 , Final_F1_89 , Final_F1_91 , Final_F1_93 , Final_F1_95
, Final_F1_121 , Final_F1_123 , Final_F1_125 , Final_F1_127 , Final_F1_129 , Final_F1_131 , Final_F1_133 , Final_F1_135 , Final_F1_137 , Final_F1_139 , Final_F1_141 , Final_F1_143
, Final_F1_169 , Final_F1_171 , Final_F1_173 , Final_F1_175 , Final_F1_177 , Final_F1_179 , Final_F1_181 , Final_F1_183 , Final_F1_185 , Final_F1_187 , Final_F1_189 , Final_F1_191
, Final_F1_217 , Final_F1_219 , Final_F1_221 , Final_F1_223 , Final_F1_225 , Final_F1_227 , Final_F1_229 , Final_F1_231 , Final_F1_233 , Final_F1_235 , Final_F1_237 , Final_F1_239
, Final_F1_265 , Final_F1_267 , Final_F1_269 , Final_F1_271 , Final_F1_273 , Final_F1_275 , Final_F1_277 , Final_F1_279 , Final_F1_281 , Final_F1_283 , Final_F1_285 , Final_F1_287
, Final_F1_313 , Final_F1_315 , Final_F1_317 , Final_F1_319 , Final_F1_321 , Final_F1_323 , Final_F1_325 , Final_F1_327 , Final_F1_329 , Final_F1_331 , Final_F1_333 , Final_F1_335
, Final_F1_361 , Final_F1_363 , Final_F1_365 , Final_F1_367 , Final_F1_369 , Final_F1_371 , Final_F1_373 , Final_F1_375 , Final_F1_377 , Final_F1_379 , Final_F1_381 , Final_F1_383
, Final_F1_409 , Final_F1_411 , Final_F1_413 , Final_F1_415 , Final_F1_417 , Final_F1_419 , Final_F1_421 , Final_F1_423 , Final_F1_425 , Final_F1_427 , Final_F1_429 , Final_F1_431
, Final_F1_457 , Final_F1_459 , Final_F1_461 , Final_F1_463 , Final_F1_465 , Final_F1_467 , Final_F1_469 , Final_F1_471 , Final_F1_473 , Final_F1_475 , Final_F1_477 , Final_F1_479
, Final_F1_505 , Final_F1_507 , Final_F1_509 , Final_F1_511 , Final_F1_513 , Final_F1_515 , Final_F1_517 , Final_F1_519 , Final_F1_521 , Final_F1_523 , Final_F1_525 , Final_F1_527
, Final_F1_553 , Final_F1_555 , Final_F1_557 , Final_F1_559 , Final_F1_561 , Final_F1_563 , Final_F1_565 , Final_F1_567 , Final_F1_569 , Final_F1_571 , Final_F1_573 , Final_F1_575
, superADDRESS, SuperMuxOut_F1_4);
*/


//COMPARATOR_MAX_TRY F1_1_1 (clk, SuperMuxOut_F1_1, SuperMuxOut_F1_2, SuperMuxOut_F1_3, SuperMuxOut_F1_4 , CompOut_F1 );
COMPARATOR_MAX_TRY_tssssst F1_1_1 (clk, RELUout_F1_1_1, RELUout_F1_1_2, RELUout_F1_2_1, RELUout_F1_2_2 , CompOut_F1 );
////
/*

SUPERMUXMODULE_MAXPOOL1_2by2_340 F2_1_1_1 
( Final_F2_0 , Final_F2_2 , Final_F2_4 , Final_F2_6 , Final_F2_8 , Final_F2_10 , Final_F2_12 , Final_F2_14 , Final_F2_16 , Final_F2_18 , Final_F2_20 , Final_F2_22
, Final_F2_48 , Final_F2_50 , Final_F2_52 , Final_F2_54 , Final_F2_56 , Final_F2_58 , Final_F2_60 , Final_F2_62 , Final_F2_64 , Final_F2_66 , Final_F2_68 , Final_F2_70
, Final_F2_96 , Final_F2_98 , Final_F2_100 , Final_F2_102 , Final_F2_104 , Final_F2_106 , Final_F2_108 , Final_F2_110 , Final_F2_112 , Final_F2_114 , Final_F2_116 , Final_F2_118
, Final_F2_144 , Final_F2_146 , Final_F2_148 , Final_F2_150 , Final_F2_152 , Final_F2_154 , Final_F2_156 , Final_F2_158 , Final_F2_160 , Final_F2_162 , Final_F2_164 , Final_F2_166
, Final_F2_192 , Final_F2_194 , Final_F2_196 , Final_F2_198 , Final_F2_200 , Final_F2_202 , Final_F2_204 , Final_F2_206 , Final_F2_208 , Final_F2_210 , Final_F2_212 , Final_F2_214
, Final_F2_240 , Final_F2_242 , Final_F2_244 , Final_F2_246 , Final_F2_248 , Final_F2_250 , Final_F2_252 , Final_F2_254 , Final_F2_256 , Final_F2_258 , Final_F2_260 , Final_F2_262
, Final_F2_288 , Final_F2_290 , Final_F2_292 , Final_F2_294 , Final_F2_296 , Final_F2_298 , Final_F2_300 , Final_F2_302 , Final_F2_304 , Final_F2_306 , Final_F2_308 , Final_F2_310
, Final_F2_336 , Final_F2_338 , Final_F2_340 , Final_F2_342 , Final_F2_344 , Final_F2_346 , Final_F2_348 , Final_F2_350 , Final_F2_352 , Final_F2_354 , Final_F2_356 , Final_F2_358
, Final_F2_384 , Final_F2_386 , Final_F2_388 , Final_F2_390 , Final_F2_392 , Final_F2_394 , Final_F2_396 , Final_F2_398 , Final_F2_400 , Final_F2_402 , Final_F2_404 , Final_F2_406
, Final_F2_432 , Final_F2_434 , Final_F2_436 , Final_F2_438 , Final_F2_440 , Final_F2_442 , Final_F2_444 , Final_F2_446 , Final_F2_448 , Final_F2_450 , Final_F2_452 , Final_F2_454
, Final_F2_480 , Final_F2_482 , Final_F2_484 , Final_F2_486 , Final_F2_488 , Final_F2_490 , Final_F2_492 , Final_F2_494 , Final_F2_496 , Final_F2_498 , Final_F2_500 , Final_F2_502
, Final_F2_528 , Final_F2_530 , Final_F2_532 , Final_F2_534 , Final_F2_536 , Final_F2_538 , Final_F2_540 , Final_F2_542 , Final_F2_544 , Final_F2_546 , Final_F2_548 , Final_F2_550
, superADDRESS, SuperMuxOut_F2_1);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F2_1_1_2 
( Final_F2_1 , Final_F2_3 , Final_F2_5 , Final_F2_7 , Final_F2_9 , Final_F2_11 , Final_F2_13 , Final_F2_15 , Final_F2_17 , Final_F2_19 , Final_F2_21 , Final_F2_23
, Final_F2_49 , Final_F2_51 , Final_F2_53 , Final_F2_55 , Final_F2_57 , Final_F2_59 , Final_F2_61 , Final_F2_63 , Final_F2_65 , Final_F2_67 , Final_F2_69 , Final_F2_71
, Final_F2_97 , Final_F2_99 , Final_F2_101 , Final_F2_103 , Final_F2_105 , Final_F2_107 , Final_F2_109 , Final_F2_111 , Final_F2_113 , Final_F2_115 , Final_F2_117 , Final_F2_119
, Final_F2_145 , Final_F2_147 , Final_F2_149 , Final_F2_151 , Final_F2_153 , Final_F2_155 , Final_F2_157 , Final_F2_159 , Final_F2_161 , Final_F2_163 , Final_F2_165 , Final_F2_167
, Final_F2_193 , Final_F2_195 , Final_F2_197 , Final_F2_199 , Final_F2_201 , Final_F2_203 , Final_F2_205 , Final_F2_207 , Final_F2_209 , Final_F2_211 , Final_F2_213 , Final_F2_215
, Final_F2_241 , Final_F2_243 , Final_F2_245 , Final_F2_247 , Final_F2_249 , Final_F2_251 , Final_F2_253 , Final_F2_255 , Final_F2_257 , Final_F2_259 , Final_F2_261 , Final_F2_263
, Final_F2_289 , Final_F2_291 , Final_F2_293 , Final_F2_295 , Final_F2_297 , Final_F2_299 , Final_F2_301 , Final_F2_303 , Final_F2_305 , Final_F2_307 , Final_F2_309 , Final_F2_311
, Final_F2_337 , Final_F2_339 , Final_F2_341 , Final_F2_343 , Final_F2_345 , Final_F2_347 , Final_F2_349 , Final_F2_351 , Final_F2_353 , Final_F2_355 , Final_F2_357 , Final_F2_359
, Final_F2_385 , Final_F2_387 , Final_F2_389 , Final_F2_391 , Final_F2_393 , Final_F2_395 , Final_F2_397 , Final_F2_399 , Final_F2_401 , Final_F2_403 , Final_F2_405 , Final_F2_407
, Final_F2_433 , Final_F2_435 , Final_F2_437 , Final_F2_439 , Final_F2_441 , Final_F2_443 , Final_F2_445 , Final_F2_447 , Final_F2_449 , Final_F2_451 , Final_F2_453 , Final_F2_455
, Final_F2_481 , Final_F2_483 , Final_F2_485 , Final_F2_487 , Final_F2_489 , Final_F2_491 , Final_F2_493 , Final_F2_495 , Final_F2_497 , Final_F2_499 , Final_F2_501 , Final_F2_503
, Final_F2_529 , Final_F2_531 , Final_F2_533 , Final_F2_535 , Final_F2_537 , Final_F2_539 , Final_F2_541 , Final_F2_543 , Final_F2_545 , Final_F2_547 , Final_F2_549 , Final_F2_551
, superADDRESS, SuperMuxOut_F2_2);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F2_1_1_3 
( Final_F2_24 , Final_F2_26 , Final_F2_28 , Final_F2_30 , Final_F2_32 , Final_F2_34 , Final_F2_36 , Final_F2_38 , Final_F2_40 , Final_F2_42 , Final_F2_44 , Final_F2_46
, Final_F2_72 , Final_F2_74 , Final_F2_76 , Final_F2_78 , Final_F2_80 , Final_F2_82 , Final_F2_84 , Final_F2_86 , Final_F2_88 , Final_F2_90 , Final_F2_92 , Final_F2_94
, Final_F2_120 , Final_F2_122 , Final_F2_124 , Final_F2_126 , Final_F2_128 , Final_F2_130 , Final_F2_132 , Final_F2_134 , Final_F2_136 , Final_F2_138 , Final_F2_140 , Final_F2_142
, Final_F2_168 , Final_F2_170 , Final_F2_172 , Final_F2_174 , Final_F2_176 , Final_F2_178 , Final_F2_180 , Final_F2_182 , Final_F2_184 , Final_F2_186 , Final_F2_188 , Final_F2_190
, Final_F2_216 , Final_F2_218 , Final_F2_220 , Final_F2_222 , Final_F2_224 , Final_F2_226 , Final_F2_228 , Final_F2_230 , Final_F2_232 , Final_F2_234 , Final_F2_236 , Final_F2_238
, Final_F2_264 , Final_F2_266 , Final_F2_268 , Final_F2_270 , Final_F2_272 , Final_F2_274 , Final_F2_276 , Final_F2_278 , Final_F2_280 , Final_F2_282 , Final_F2_284 , Final_F2_286
, Final_F2_312 , Final_F2_314 , Final_F2_316 , Final_F2_318 , Final_F2_320 , Final_F2_322 , Final_F2_324 , Final_F2_326 , Final_F2_328 , Final_F2_330 , Final_F2_332 , Final_F2_334
, Final_F2_360 , Final_F2_362 , Final_F2_364 , Final_F2_366 , Final_F2_368 , Final_F2_370 , Final_F2_372 , Final_F2_374 , Final_F2_376 , Final_F2_378 , Final_F2_380 , Final_F2_382
, Final_F2_408 , Final_F2_410 , Final_F2_412 , Final_F2_414 , Final_F2_416 , Final_F2_418 , Final_F2_420 , Final_F2_422 , Final_F2_424 , Final_F2_426 , Final_F2_428 , Final_F2_430
, Final_F2_456 , Final_F2_458 , Final_F2_460 , Final_F2_462 , Final_F2_464 , Final_F2_466 , Final_F2_468 , Final_F2_470 , Final_F2_472 , Final_F2_474 , Final_F2_476 , Final_F2_478
, Final_F2_504 , Final_F2_506 , Final_F2_508 , Final_F2_510 , Final_F2_512 , Final_F2_514 , Final_F2_516 , Final_F2_518 , Final_F2_520 , Final_F2_522 , Final_F2_524 , Final_F2_526
, Final_F2_552 , Final_F2_554 , Final_F2_556 , Final_F2_558 , Final_F2_560 , Final_F2_562 , Final_F2_564 , Final_F2_566 , Final_F2_568 , Final_F2_570 , Final_F2_572 , Final_F2_574
, superADDRESS, SuperMuxOut_F2_3);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F2_1_1_4
( Final_F2_25 , Final_F2_27 , Final_F2_29 , Final_F2_31 , Final_F2_33 , Final_F2_35 , Final_F2_37 , Final_F2_39 , Final_F2_41 , Final_F2_43 , Final_F2_45 , Final_F2_47
, Final_F2_73 , Final_F2_75 , Final_F2_77 , Final_F2_79 , Final_F2_81 , Final_F2_83 , Final_F2_85 , Final_F2_87 , Final_F2_89 , Final_F2_91 , Final_F2_93 , Final_F2_95
, Final_F2_121 , Final_F2_123 , Final_F2_125 , Final_F2_127 , Final_F2_129 , Final_F2_131 , Final_F2_133 , Final_F2_135 , Final_F2_137 , Final_F2_139 , Final_F2_141 , Final_F2_143
, Final_F2_169 , Final_F2_171 , Final_F2_173 , Final_F2_175 , Final_F2_177 , Final_F2_179 , Final_F2_181 , Final_F2_183 , Final_F2_185 , Final_F2_187 , Final_F2_189 , Final_F2_191
, Final_F2_217 , Final_F2_219 , Final_F2_221 , Final_F2_223 , Final_F2_225 , Final_F2_227 , Final_F2_229 , Final_F2_231 , Final_F2_233 , Final_F2_235 , Final_F2_237 , Final_F2_239
, Final_F2_265 , Final_F2_267 , Final_F2_269 , Final_F2_271 , Final_F2_273 , Final_F2_275 , Final_F2_277 , Final_F2_279 , Final_F2_281 , Final_F2_283 , Final_F2_285 , Final_F2_287
, Final_F2_313 , Final_F2_315 , Final_F2_317 , Final_F2_319 , Final_F2_321 , Final_F2_323 , Final_F2_325 , Final_F2_327 , Final_F2_329 , Final_F2_331 , Final_F2_333 , Final_F2_335
, Final_F2_361 , Final_F2_363 , Final_F2_365 , Final_F2_367 , Final_F2_369 , Final_F2_371 , Final_F2_373 , Final_F2_375 , Final_F2_377 , Final_F2_379 , Final_F2_381 , Final_F2_383
, Final_F2_409 , Final_F2_411 , Final_F2_413 , Final_F2_415 , Final_F2_417 , Final_F2_419 , Final_F2_421 , Final_F2_423 , Final_F2_425 , Final_F2_427 , Final_F2_429 , Final_F2_431
, Final_F2_457 , Final_F2_459 , Final_F2_461 , Final_F2_463 , Final_F2_465 , Final_F2_467 , Final_F2_469 , Final_F2_471 , Final_F2_473 , Final_F2_475 , Final_F2_477 , Final_F2_479
, Final_F2_505 , Final_F2_507 , Final_F2_509 , Final_F2_511 , Final_F2_513 , Final_F2_515 , Final_F2_517 , Final_F2_519 , Final_F2_521 , Final_F2_523 , Final_F2_525 , Final_F2_527
, Final_F2_553 , Final_F2_555 , Final_F2_557 , Final_F2_559 , Final_F2_561 , Final_F2_563 , Final_F2_565 , Final_F2_567 , Final_F2_569 , Final_F2_571 , Final_F2_573 , Final_F2_575
, superADDRESS, SuperMuxOut_F2_4);

*/
//COMPARATOR_MAX_TRY F2_1_1 (clk, SuperMuxOut_F2_1, SuperMuxOut_F2_2, SuperMuxOut_F2_3, SuperMuxOut_F2_4 , CompOut_F2 );
COMPARATOR_MAX_TRY_tssssst F2_1_1 (clk, RELUout_F2_1_1, RELUout_F2_1_2, RELUout_F2_2_1, RELUout_F2_2_2 , CompOut_F2 );

///
/*
SUPERMUXMODULE_MAXPOOL1_2by2_340 F3_1_1_1 
( Final_F3_0 , Final_F3_2 , Final_F3_4 , Final_F3_6 , Final_F3_8 , Final_F3_10 , Final_F3_12 , Final_F3_14 , Final_F3_16 , Final_F3_18 , Final_F3_20 , Final_F3_22
, Final_F3_48 , Final_F3_50 , Final_F3_52 , Final_F3_54 , Final_F3_56 , Final_F3_58 , Final_F3_60 , Final_F3_62 , Final_F3_64 , Final_F3_66 , Final_F3_68 , Final_F3_70
, Final_F3_96 , Final_F3_98 , Final_F3_100 , Final_F3_102 , Final_F3_104 , Final_F3_106 , Final_F3_108 , Final_F3_110 , Final_F3_112 , Final_F3_114 , Final_F3_116 , Final_F3_118
, Final_F3_144 , Final_F3_146 , Final_F3_148 , Final_F3_150 , Final_F3_152 , Final_F3_154 , Final_F3_156 , Final_F3_158 , Final_F3_160 , Final_F3_162 , Final_F3_164 , Final_F3_166
, Final_F3_192 , Final_F3_194 , Final_F3_196 , Final_F3_198 , Final_F3_200 , Final_F3_202 , Final_F3_204 , Final_F3_206 , Final_F3_208 , Final_F3_210 , Final_F3_212 , Final_F3_214
, Final_F3_240 , Final_F3_242 , Final_F3_244 , Final_F3_246 , Final_F3_248 , Final_F3_250 , Final_F3_252 , Final_F3_254 , Final_F3_256 , Final_F3_258 , Final_F3_260 , Final_F3_262
, Final_F3_288 , Final_F3_290 , Final_F3_292 , Final_F3_294 , Final_F3_296 , Final_F3_298 , Final_F3_300 , Final_F3_302 , Final_F3_304 , Final_F3_306 , Final_F3_308 , Final_F3_310
, Final_F3_336 , Final_F3_338 , Final_F3_340 , Final_F3_342 , Final_F3_344 , Final_F3_346 , Final_F3_348 , Final_F3_350 , Final_F3_352 , Final_F3_354 , Final_F3_356 , Final_F3_358
, Final_F3_384 , Final_F3_386 , Final_F3_388 , Final_F3_390 , Final_F3_392 , Final_F3_394 , Final_F3_396 , Final_F3_398 , Final_F3_400 , Final_F3_402 , Final_F3_404 , Final_F3_406
, Final_F3_432 , Final_F3_434 , Final_F3_436 , Final_F3_438 , Final_F3_440 , Final_F3_442 , Final_F3_444 , Final_F3_446 , Final_F3_448 , Final_F3_450 , Final_F3_452 , Final_F3_454
, Final_F3_480 , Final_F3_482 , Final_F3_484 , Final_F3_486 , Final_F3_488 , Final_F3_490 , Final_F3_492 , Final_F3_494 , Final_F3_496 , Final_F3_498 , Final_F3_500 , Final_F3_502
, Final_F3_528 , Final_F3_530 , Final_F3_532 , Final_F3_534 , Final_F3_536 , Final_F3_538 , Final_F3_540 , Final_F3_542 , Final_F3_544 , Final_F3_546 , Final_F3_548 , Final_F3_550
, superADDRESS, SuperMuxOut_F3_1);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F3_1_1_2 
( Final_F3_1 , Final_F3_3 , Final_F3_5 , Final_F3_7 , Final_F3_9 , Final_F3_11 , Final_F3_13 , Final_F3_15 , Final_F3_17 , Final_F3_19 , Final_F3_21 , Final_F3_23
, Final_F3_49 , Final_F3_51 , Final_F3_53 , Final_F3_55 , Final_F3_57 , Final_F3_59 , Final_F3_61 , Final_F3_63 , Final_F3_65 , Final_F3_67 , Final_F3_69 , Final_F3_71
, Final_F3_97 , Final_F3_99 , Final_F3_101 , Final_F3_103 , Final_F3_105 , Final_F3_107 , Final_F3_109 , Final_F3_111 , Final_F3_113 , Final_F3_115 , Final_F3_117 , Final_F3_119
, Final_F3_145 , Final_F3_147 , Final_F3_149 , Final_F3_151 , Final_F3_153 , Final_F3_155 , Final_F3_157 , Final_F3_159 , Final_F3_161 , Final_F3_163 , Final_F3_165 , Final_F3_167
, Final_F3_193 , Final_F3_195 , Final_F3_197 , Final_F3_199 , Final_F3_201 , Final_F3_203 , Final_F3_205 , Final_F3_207 , Final_F3_209 , Final_F3_211 , Final_F3_213 , Final_F3_215
, Final_F3_241 , Final_F3_243 , Final_F3_245 , Final_F3_247 , Final_F3_249 , Final_F3_251 , Final_F3_253 , Final_F3_255 , Final_F3_257 , Final_F3_259 , Final_F3_261 , Final_F3_263
, Final_F3_289 , Final_F3_291 , Final_F3_293 , Final_F3_295 , Final_F3_297 , Final_F3_299 , Final_F3_301 , Final_F3_303 , Final_F3_305 , Final_F3_307 , Final_F3_309 , Final_F3_311
, Final_F3_337 , Final_F3_339 , Final_F3_341 , Final_F3_343 , Final_F3_345 , Final_F3_347 , Final_F3_349 , Final_F3_351 , Final_F3_353 , Final_F3_355 , Final_F3_357 , Final_F3_359
, Final_F3_385 , Final_F3_387 , Final_F3_389 , Final_F3_391 , Final_F3_393 , Final_F3_395 , Final_F3_397 , Final_F3_399 , Final_F3_401 , Final_F3_403 , Final_F3_405 , Final_F3_407
, Final_F3_433 , Final_F3_435 , Final_F3_437 , Final_F3_439 , Final_F3_441 , Final_F3_443 , Final_F3_445 , Final_F3_447 , Final_F3_449 , Final_F3_451 , Final_F3_453 , Final_F3_455
, Final_F3_481 , Final_F3_483 , Final_F3_485 , Final_F3_487 , Final_F3_489 , Final_F3_491 , Final_F3_493 , Final_F3_495 , Final_F3_497 , Final_F3_499 , Final_F3_501 , Final_F3_503
, Final_F3_529 , Final_F3_531 , Final_F3_533 , Final_F3_535 , Final_F3_537 , Final_F3_539 , Final_F3_541 , Final_F3_543 , Final_F3_545 , Final_F3_547 , Final_F3_549 , Final_F3_551
, superADDRESS, SuperMuxOut_F3_2);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F3_1_1_3 
( Final_F3_24 , Final_F3_26 , Final_F3_28 , Final_F3_30 , Final_F3_32 , Final_F3_34 , Final_F3_36 , Final_F3_38 , Final_F3_40 , Final_F3_42 , Final_F3_44 , Final_F3_46
, Final_F3_72 , Final_F3_74 , Final_F3_76 , Final_F3_78 , Final_F3_80 , Final_F3_82 , Final_F3_84 , Final_F3_86 , Final_F3_88 , Final_F3_90 , Final_F3_92 , Final_F3_94
, Final_F3_120 , Final_F3_122 , Final_F3_124 , Final_F3_126 , Final_F3_128 , Final_F3_130 , Final_F3_132 , Final_F3_134 , Final_F3_136 , Final_F3_138 , Final_F3_140 , Final_F3_142
, Final_F3_168 , Final_F3_170 , Final_F3_172 , Final_F3_174 , Final_F3_176 , Final_F3_178 , Final_F3_180 , Final_F3_182 , Final_F3_184 , Final_F3_186 , Final_F3_188 , Final_F3_190
, Final_F3_216 , Final_F3_218 , Final_F3_220 , Final_F3_222 , Final_F3_224 , Final_F3_226 , Final_F3_228 , Final_F3_230 , Final_F3_232 , Final_F3_234 , Final_F3_236 , Final_F3_238
, Final_F3_264 , Final_F3_266 , Final_F3_268 , Final_F3_270 , Final_F3_272 , Final_F3_274 , Final_F3_276 , Final_F3_278 , Final_F3_280 , Final_F3_282 , Final_F3_284 , Final_F3_286
, Final_F3_312 , Final_F3_314 , Final_F3_316 , Final_F3_318 , Final_F3_320 , Final_F3_322 , Final_F3_324 , Final_F3_326 , Final_F3_328 , Final_F3_330 , Final_F3_332 , Final_F3_334
, Final_F3_360 , Final_F3_362 , Final_F3_364 , Final_F3_366 , Final_F3_368 , Final_F3_370 , Final_F3_372 , Final_F3_374 , Final_F3_376 , Final_F3_378 , Final_F3_380 , Final_F3_382
, Final_F3_408 , Final_F3_410 , Final_F3_412 , Final_F3_414 , Final_F3_416 , Final_F3_418 , Final_F3_420 , Final_F3_422 , Final_F3_424 , Final_F3_426 , Final_F3_428 , Final_F3_430
, Final_F3_456 , Final_F3_458 , Final_F3_460 , Final_F3_462 , Final_F3_464 , Final_F3_466 , Final_F3_468 , Final_F3_470 , Final_F3_472 , Final_F3_474 , Final_F3_476 , Final_F3_478
, Final_F3_504 , Final_F3_506 , Final_F3_508 , Final_F3_510 , Final_F3_512 , Final_F3_514 , Final_F3_516 , Final_F3_518 , Final_F3_520 , Final_F3_522 , Final_F3_524 , Final_F3_526
, Final_F3_552 , Final_F3_554 , Final_F3_556 , Final_F3_558 , Final_F3_560 , Final_F3_562 , Final_F3_564 , Final_F3_566 , Final_F3_568 , Final_F3_570 , Final_F3_572 , Final_F3_574
, superADDRESS, SuperMuxOut_F3_3);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F3_1_1_4
( Final_F3_25 , Final_F3_27 , Final_F3_29 , Final_F3_31 , Final_F3_33 , Final_F3_35 , Final_F3_37 , Final_F3_39 , Final_F3_41 , Final_F3_43 , Final_F3_45 , Final_F3_47
, Final_F3_73 , Final_F3_75 , Final_F3_77 , Final_F3_79 , Final_F3_81 , Final_F3_83 , Final_F3_85 , Final_F3_87 , Final_F3_89 , Final_F3_91 , Final_F3_93 , Final_F3_95
, Final_F3_121 , Final_F3_123 , Final_F3_125 , Final_F3_127 , Final_F3_129 , Final_F3_131 , Final_F3_133 , Final_F3_135 , Final_F3_137 , Final_F3_139 , Final_F3_141 , Final_F3_143
, Final_F3_169 , Final_F3_171 , Final_F3_173 , Final_F3_175 , Final_F3_177 , Final_F3_179 , Final_F3_181 , Final_F3_183 , Final_F3_185 , Final_F3_187 , Final_F3_189 , Final_F3_191
, Final_F3_217 , Final_F3_219 , Final_F3_221 , Final_F3_223 , Final_F3_225 , Final_F3_227 , Final_F3_229 , Final_F3_231 , Final_F3_233 , Final_F3_235 , Final_F3_237 , Final_F3_239
, Final_F3_265 , Final_F3_267 , Final_F3_269 , Final_F3_271 , Final_F3_273 , Final_F3_275 , Final_F3_277 , Final_F3_279 , Final_F3_281 , Final_F3_283 , Final_F3_285 , Final_F3_287
, Final_F3_313 , Final_F3_315 , Final_F3_317 , Final_F3_319 , Final_F3_321 , Final_F3_323 , Final_F3_325 , Final_F3_327 , Final_F3_329 , Final_F3_331 , Final_F3_333 , Final_F3_335
, Final_F3_361 , Final_F3_363 , Final_F3_365 , Final_F3_367 , Final_F3_369 , Final_F3_371 , Final_F3_373 , Final_F3_375 , Final_F3_377 , Final_F3_379 , Final_F3_381 , Final_F3_383
, Final_F3_409 , Final_F3_411 , Final_F3_413 , Final_F3_415 , Final_F3_417 , Final_F3_419 , Final_F3_421 , Final_F3_423 , Final_F3_425 , Final_F3_427 , Final_F3_429 , Final_F3_431
, Final_F3_457 , Final_F3_459 , Final_F3_461 , Final_F3_463 , Final_F3_465 , Final_F3_467 , Final_F3_469 , Final_F3_471 , Final_F3_473 , Final_F3_475 , Final_F3_477 , Final_F3_479
, Final_F3_505 , Final_F3_507 , Final_F3_509 , Final_F3_511 , Final_F3_513 , Final_F3_515 , Final_F3_517 , Final_F3_519 , Final_F3_521 , Final_F3_523 , Final_F3_525 , Final_F3_527
, Final_F3_553 , Final_F3_555 , Final_F3_557 , Final_F3_559 , Final_F3_561 , Final_F3_563 , Final_F3_565 , Final_F3_567 , Final_F3_569 , Final_F3_571 , Final_F3_573 , Final_F3_575
, superADDRESS, SuperMuxOut_F3_4);
*/

//COMPARATOR_MAX_TRY F3_1_1 (clk, SuperMuxOut_F3_1, SuperMuxOut_F3_2, SuperMuxOut_F3_3, SuperMuxOut_F3_4 , CompOut_F3 );
COMPARATOR_MAX_TRY_tssssst F3_1_1 (clk, RELUout_F3_1_1, RELUout_F3_1_2, RELUout_F3_2_1, RELUout_F3_2_2 , CompOut_F3 );
////
/*
SUPERMUXMODULE_MAXPOOL1_2by2_340 F4_1_1_1 
( Final_F4_0 , Final_F4_2 , Final_F4_4 , Final_F4_6 , Final_F4_8 , Final_F4_10 , Final_F4_12 , Final_F4_14 , Final_F4_16 , Final_F4_18 , Final_F4_20 , Final_F4_22
, Final_F4_48 , Final_F4_50 , Final_F4_52 , Final_F4_54 , Final_F4_56 , Final_F4_58 , Final_F4_60 , Final_F4_62 , Final_F4_64 , Final_F4_66 , Final_F4_68 , Final_F4_70
, Final_F4_96 , Final_F4_98 , Final_F4_100 , Final_F4_102 , Final_F4_104 , Final_F4_106 , Final_F4_108 , Final_F4_110 , Final_F4_112 , Final_F4_114 , Final_F4_116 , Final_F4_118
, Final_F4_144 , Final_F4_146 , Final_F4_148 , Final_F4_150 , Final_F4_152 , Final_F4_154 , Final_F4_156 , Final_F4_158 , Final_F4_160 , Final_F4_162 , Final_F4_164 , Final_F4_166
, Final_F4_192 , Final_F4_194 , Final_F4_196 , Final_F4_198 , Final_F4_200 , Final_F4_202 , Final_F4_204 , Final_F4_206 , Final_F4_208 , Final_F4_210 , Final_F4_212 , Final_F4_214
, Final_F4_240 , Final_F4_242 , Final_F4_244 , Final_F4_246 , Final_F4_248 , Final_F4_250 , Final_F4_252 , Final_F4_254 , Final_F4_256 , Final_F4_258 , Final_F4_260 , Final_F4_262
, Final_F4_288 , Final_F4_290 , Final_F4_292 , Final_F4_294 , Final_F4_296 , Final_F4_298 , Final_F4_300 , Final_F4_302 , Final_F4_304 , Final_F4_306 , Final_F4_308 , Final_F4_310
, Final_F4_336 , Final_F4_338 , Final_F4_340 , Final_F4_342 , Final_F4_344 , Final_F4_346 , Final_F4_348 , Final_F4_350 , Final_F4_352 , Final_F4_354 , Final_F4_356 , Final_F4_358
, Final_F4_384 , Final_F4_386 , Final_F4_388 , Final_F4_390 , Final_F4_392 , Final_F4_394 , Final_F4_396 , Final_F4_398 , Final_F4_400 , Final_F4_402 , Final_F4_404 , Final_F4_406
, Final_F4_432 , Final_F4_434 , Final_F4_436 , Final_F4_438 , Final_F4_440 , Final_F4_442 , Final_F4_444 , Final_F4_446 , Final_F4_448 , Final_F4_450 , Final_F4_452 , Final_F4_454
, Final_F4_480 , Final_F4_482 , Final_F4_484 , Final_F4_486 , Final_F4_488 , Final_F4_490 , Final_F4_492 , Final_F4_494 , Final_F4_496 , Final_F4_498 , Final_F4_500 , Final_F4_502
, Final_F4_528 , Final_F4_530 , Final_F4_532 , Final_F4_534 , Final_F4_536 , Final_F4_538 , Final_F4_540 , Final_F4_542 , Final_F4_544 , Final_F4_546 , Final_F4_548 , Final_F4_550
, superADDRESS, SuperMuxOut_F4_1);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F4_1_1_2 
( Final_F4_1 , Final_F4_3 , Final_F4_5 , Final_F4_7 , Final_F4_9 , Final_F4_11 , Final_F4_13 , Final_F4_15 , Final_F4_17 , Final_F4_19 , Final_F4_21 , Final_F4_23
, Final_F4_49 , Final_F4_51 , Final_F4_53 , Final_F4_55 , Final_F4_57 , Final_F4_59 , Final_F4_61 , Final_F4_63 , Final_F4_65 , Final_F4_67 , Final_F4_69 , Final_F4_71
, Final_F4_97 , Final_F4_99 , Final_F4_101 , Final_F4_103 , Final_F4_105 , Final_F4_107 , Final_F4_109 , Final_F4_111 , Final_F4_113 , Final_F4_115 , Final_F4_117 , Final_F4_119
, Final_F4_145 , Final_F4_147 , Final_F4_149 , Final_F4_151 , Final_F4_153 , Final_F4_155 , Final_F4_157 , Final_F4_159 , Final_F4_161 , Final_F4_163 , Final_F4_165 , Final_F4_167
, Final_F4_193 , Final_F4_195 , Final_F4_197 , Final_F4_199 , Final_F4_201 , Final_F4_203 , Final_F4_205 , Final_F4_207 , Final_F4_209 , Final_F4_211 , Final_F4_213 , Final_F4_215
, Final_F4_241 , Final_F4_243 , Final_F4_245 , Final_F4_247 , Final_F4_249 , Final_F4_251 , Final_F4_253 , Final_F4_255 , Final_F4_257 , Final_F4_259 , Final_F4_261 , Final_F4_263
, Final_F4_289 , Final_F4_291 , Final_F4_293 , Final_F4_295 , Final_F4_297 , Final_F4_299 , Final_F4_301 , Final_F4_303 , Final_F4_305 , Final_F4_307 , Final_F4_309 , Final_F4_311
, Final_F4_337 , Final_F4_339 , Final_F4_341 , Final_F4_343 , Final_F4_345 , Final_F4_347 , Final_F4_349 , Final_F4_351 , Final_F4_353 , Final_F4_355 , Final_F4_357 , Final_F4_359
, Final_F4_385 , Final_F4_387 , Final_F4_389 , Final_F4_391 , Final_F4_393 , Final_F4_395 , Final_F4_397 , Final_F4_399 , Final_F4_401 , Final_F4_403 , Final_F4_405 , Final_F4_407
, Final_F4_433 , Final_F4_435 , Final_F4_437 , Final_F4_439 , Final_F4_441 , Final_F4_443 , Final_F4_445 , Final_F4_447 , Final_F4_449 , Final_F4_451 , Final_F4_453 , Final_F4_455
, Final_F4_481 , Final_F4_483 , Final_F4_485 , Final_F4_487 , Final_F4_489 , Final_F4_491 , Final_F4_493 , Final_F4_495 , Final_F4_497 , Final_F4_499 , Final_F4_501 , Final_F4_503
, Final_F4_529 , Final_F4_531 , Final_F4_533 , Final_F4_535 , Final_F4_537 , Final_F4_539 , Final_F4_541 , Final_F4_543 , Final_F4_545 , Final_F4_547 , Final_F4_549 , Final_F4_551
, superADDRESS, SuperMuxOut_F4_2);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F4_1_1_3 
( Final_F4_24 , Final_F4_26 , Final_F4_28 , Final_F4_30 , Final_F4_32 , Final_F4_34 , Final_F4_36 , Final_F4_38 , Final_F4_40 , Final_F4_42 , Final_F4_44 , Final_F4_46
, Final_F4_72 , Final_F4_74 , Final_F4_76 , Final_F4_78 , Final_F4_80 , Final_F4_82 , Final_F4_84 , Final_F4_86 , Final_F4_88 , Final_F4_90 , Final_F4_92 , Final_F4_94
, Final_F4_120 , Final_F4_122 , Final_F4_124 , Final_F4_126 , Final_F4_128 , Final_F4_130 , Final_F4_132 , Final_F4_134 , Final_F4_136 , Final_F4_138 , Final_F4_140 , Final_F4_142
, Final_F4_168 , Final_F4_170 , Final_F4_172 , Final_F4_174 , Final_F4_176 , Final_F4_178 , Final_F4_180 , Final_F4_182 , Final_F4_184 , Final_F4_186 , Final_F4_188 , Final_F4_190
, Final_F4_216 , Final_F4_218 , Final_F4_220 , Final_F4_222 , Final_F4_224 , Final_F4_226 , Final_F4_228 , Final_F4_230 , Final_F4_232 , Final_F4_234 , Final_F4_236 , Final_F4_238
, Final_F4_264 , Final_F4_266 , Final_F4_268 , Final_F4_270 , Final_F4_272 , Final_F4_274 , Final_F4_276 , Final_F4_278 , Final_F4_280 , Final_F4_282 , Final_F4_284 , Final_F4_286
, Final_F4_312 , Final_F4_314 , Final_F4_316 , Final_F4_318 , Final_F4_320 , Final_F4_322 , Final_F4_324 , Final_F4_326 , Final_F4_328 , Final_F4_330 , Final_F4_332 , Final_F4_334
, Final_F4_360 , Final_F4_362 , Final_F4_364 , Final_F4_366 , Final_F4_368 , Final_F4_370 , Final_F4_372 , Final_F4_374 , Final_F4_376 , Final_F4_378 , Final_F4_380 , Final_F4_382
, Final_F4_408 , Final_F4_410 , Final_F4_412 , Final_F4_414 , Final_F4_416 , Final_F4_418 , Final_F4_420 , Final_F4_422 , Final_F4_424 , Final_F4_426 , Final_F4_428 , Final_F4_430
, Final_F4_456 , Final_F4_458 , Final_F4_460 , Final_F4_462 , Final_F4_464 , Final_F4_466 , Final_F4_468 , Final_F4_470 , Final_F4_472 , Final_F4_474 , Final_F4_476 , Final_F4_478
, Final_F4_504 , Final_F4_506 , Final_F4_508 , Final_F4_510 , Final_F4_512 , Final_F4_514 , Final_F4_516 , Final_F4_518 , Final_F4_520 , Final_F4_522 , Final_F4_524 , Final_F4_526
, Final_F4_552 , Final_F4_554 , Final_F4_556 , Final_F4_558 , Final_F4_560 , Final_F4_562 , Final_F4_564 , Final_F4_566 , Final_F4_568 , Final_F4_570 , Final_F4_572 , Final_F4_574
, superADDRESS, SuperMuxOut_F4_3);
SUPERMUXMODULE_MAXPOOL1_2by2_340 F4_1_1_4
( Final_F4_25 , Final_F4_27 , Final_F4_29 , Final_F4_31 , Final_F4_33 , Final_F4_35 , Final_F4_37 , Final_F4_39 , Final_F4_41 , Final_F4_43 , Final_F4_45 , Final_F4_47
, Final_F4_73 , Final_F4_75 , Final_F4_77 , Final_F4_79 , Final_F4_81 , Final_F4_83 , Final_F4_85 , Final_F4_87 , Final_F4_89 , Final_F4_91 , Final_F4_93 , Final_F4_95
, Final_F4_121 , Final_F4_123 , Final_F4_125 , Final_F4_127 , Final_F4_129 , Final_F4_131 , Final_F4_133 , Final_F4_135 , Final_F4_137 , Final_F4_139 , Final_F4_141 , Final_F4_143
, Final_F4_169 , Final_F4_171 , Final_F4_173 , Final_F4_175 , Final_F4_177 , Final_F4_179 , Final_F4_181 , Final_F4_183 , Final_F4_185 , Final_F4_187 , Final_F4_189 , Final_F4_191
, Final_F4_217 , Final_F4_219 , Final_F4_221 , Final_F4_223 , Final_F4_225 , Final_F4_227 , Final_F4_229 , Final_F4_231 , Final_F4_233 , Final_F4_235 , Final_F4_237 , Final_F4_239
, Final_F4_265 , Final_F4_267 , Final_F4_269 , Final_F4_271 , Final_F4_273 , Final_F4_275 , Final_F4_277 , Final_F4_279 , Final_F4_281 , Final_F4_283 , Final_F4_285 , Final_F4_287
, Final_F4_313 , Final_F4_315 , Final_F4_317 , Final_F4_319 , Final_F4_321 , Final_F4_323 , Final_F4_325 , Final_F4_327 , Final_F4_329 , Final_F4_331 , Final_F4_333 , Final_F4_335
, Final_F4_361 , Final_F4_363 , Final_F4_365 , Final_F4_367 , Final_F4_369 , Final_F4_371 , Final_F4_373 , Final_F4_375 , Final_F4_377 , Final_F4_379 , Final_F4_381 , Final_F4_383
, Final_F4_409 , Final_F4_411 , Final_F4_413 , Final_F4_415 , Final_F4_417 , Final_F4_419 , Final_F4_421 , Final_F4_423 , Final_F4_425 , Final_F4_427 , Final_F4_429 , Final_F4_431
, Final_F4_457 , Final_F4_459 , Final_F4_461 , Final_F4_463 , Final_F4_465 , Final_F4_467 , Final_F4_469 , Final_F4_471 , Final_F4_473 , Final_F4_475 , Final_F4_477 , Final_F4_479
, Final_F4_505 , Final_F4_507 , Final_F4_509 , Final_F4_511 , Final_F4_513 , Final_F4_515 , Final_F4_517 , Final_F4_519 , Final_F4_521 , Final_F4_523 , Final_F4_525 , Final_F4_527
, Final_F4_553 , Final_F4_555 , Final_F4_557 , Final_F4_559 , Final_F4_561 , Final_F4_563 , Final_F4_565 , Final_F4_567 , Final_F4_569 , Final_F4_571 , Final_F4_573 , Final_F4_575
, superADDRESS, SuperMuxOut_F4_4);

*/
//COMPARATOR_MAX_TRY F4_1_1 (clk, SuperMuxOut_F4_1, SuperMuxOut_F4_2, SuperMuxOut_F4_3, SuperMuxOut_F4_4 , CompOut_F4 );
COMPARATOR_MAX_TRY_tssssst F4_1_1 (clk, RELUout_F4_1_1, RELUout_F4_1_2, RELUout_F4_2_1, RELUout_F4_2_2 , CompOut_F4 );



OneRegister MUX1_F1_RO0(clk, write2_1, CompOut_F1, REGofMAX1DataOut_F1_0 ); 
OneRegister MUX1_F1_RO1(clk, write2_2, CompOut_F1, REGofMAX1DataOut_F1_1 ); 
OneRegister MUX1_F1_RO2(clk, write2_3, CompOut_F1, REGofMAX1DataOut_F1_2 ); 
OneRegister MUX1_F1_RO3(clk, write2_4, CompOut_F1, REGofMAX1DataOut_F1_3 ); 
OneRegister MUX1_F1_RO4(clk, write2_5, CompOut_F1, REGofMAX1DataOut_F1_4 ); 
OneRegister MUX1_F1_RO5(clk, write2_6, CompOut_F1, REGofMAX1DataOut_F1_5 ); 
OneRegister MUX1_F1_RO6(clk, write2_7, CompOut_F1, REGofMAX1DataOut_F1_6 ); 
OneRegister MUX1_F1_RO7(clk, write2_8, CompOut_F1, REGofMAX1DataOut_F1_7 ); 
OneRegister MUX1_F1_RO8(clk, write2_9, CompOut_F1, REGofMAX1DataOut_F1_8 ); 
OneRegister MUX1_F1_RO9(clk, write2_10, CompOut_F1, REGofMAX1DataOut_F1_9 ); 
OneRegister MUX1_F1_RO10(clk, write2_11, CompOut_F1, REGofMAX1DataOut_F1_10 ); 
OneRegister MUX1_F1_RO11(clk, write2_12, CompOut_F1, REGofMAX1DataOut_F1_11 ); 
OneRegister MUX1_F1_RO12(clk, write2_13, CompOut_F1, REGofMAX1DataOut_F1_12 ); 
OneRegister MUX1_F1_RO13(clk, write2_14, CompOut_F1, REGofMAX1DataOut_F1_13 ); 
OneRegister MUX1_F1_RO14(clk, write2_15, CompOut_F1, REGofMAX1DataOut_F1_14 ); 
OneRegister MUX1_F1_RO15(clk, write2_16, CompOut_F1, REGofMAX1DataOut_F1_15 ); 
OneRegister MUX1_F1_RO16(clk, write2_17, CompOut_F1, REGofMAX1DataOut_F1_16 ); 
OneRegister MUX1_F1_RO17(clk, write2_18, CompOut_F1, REGofMAX1DataOut_F1_17 ); 
OneRegister MUX1_F1_RO18(clk, write2_19, CompOut_F1, REGofMAX1DataOut_F1_18 ); 
OneRegister MUX1_F1_RO19(clk, write2_20, CompOut_F1, REGofMAX1DataOut_F1_19 ); 
OneRegister MUX1_F1_RO20(clk, write2_21, CompOut_F1, REGofMAX1DataOut_F1_20 ); 
OneRegister MUX1_F1_RO21(clk, write2_22, CompOut_F1, REGofMAX1DataOut_F1_21 ); 
OneRegister MUX1_F1_RO22(clk, write2_23, CompOut_F1, REGofMAX1DataOut_F1_22 ); 
OneRegister MUX1_F1_RO23(clk, write2_24, CompOut_F1, REGofMAX1DataOut_F1_23 ); 
OneRegister MUX1_F1_RO24(clk, write2_25, CompOut_F1, REGofMAX1DataOut_F1_24 ); 
OneRegister MUX1_F1_RO25(clk, write2_26, CompOut_F1, REGofMAX1DataOut_F1_25 ); 
OneRegister MUX1_F1_RO26(clk, write2_27, CompOut_F1, REGofMAX1DataOut_F1_26 ); 
OneRegister MUX1_F1_RO27(clk, write2_28, CompOut_F1, REGofMAX1DataOut_F1_27 ); 
OneRegister MUX1_F1_RO28(clk, write2_29, CompOut_F1, REGofMAX1DataOut_F1_28 ); 
OneRegister MUX1_F1_RO29(clk, write2_30, CompOut_F1, REGofMAX1DataOut_F1_29 ); 
OneRegister MUX1_F1_RO30(clk, write2_31, CompOut_F1, REGofMAX1DataOut_F1_30 ); 
OneRegister MUX1_F1_RO31(clk, write2_32, CompOut_F1, REGofMAX1DataOut_F1_31 ); 
OneRegister MUX1_F1_RO32(clk, write2_33, CompOut_F1, REGofMAX1DataOut_F1_32 ); 
OneRegister MUX1_F1_RO33(clk, write2_34, CompOut_F1, REGofMAX1DataOut_F1_33 ); 
OneRegister MUX1_F1_RO34(clk, write2_35, CompOut_F1, REGofMAX1DataOut_F1_34 ); 
OneRegister MUX1_F1_RO35(clk, write2_36, CompOut_F1, REGofMAX1DataOut_F1_35 ); 
OneRegister MUX1_F1_RO36(clk, write2_37, CompOut_F1, REGofMAX1DataOut_F1_36 ); 
OneRegister MUX1_F1_RO37(clk, write2_38, CompOut_F1, REGofMAX1DataOut_F1_37 ); 
OneRegister MUX1_F1_RO38(clk, write2_39, CompOut_F1, REGofMAX1DataOut_F1_38 ); 
OneRegister MUX1_F1_RO39(clk, write2_40, CompOut_F1, REGofMAX1DataOut_F1_39 ); 
OneRegister MUX1_F1_RO40(clk, write2_41, CompOut_F1, REGofMAX1DataOut_F1_40 ); 
OneRegister MUX1_F1_RO41(clk, write2_42, CompOut_F1, REGofMAX1DataOut_F1_41 ); 
OneRegister MUX1_F1_RO42(clk, write2_43, CompOut_F1, REGofMAX1DataOut_F1_42 ); 
OneRegister MUX1_F1_RO43(clk, write2_44, CompOut_F1, REGofMAX1DataOut_F1_43 ); 
OneRegister MUX1_F1_RO44(clk, write2_45, CompOut_F1, REGofMAX1DataOut_F1_44 ); 
OneRegister MUX1_F1_RO45(clk, write2_46, CompOut_F1, REGofMAX1DataOut_F1_45 ); 
OneRegister MUX1_F1_RO46(clk, write2_47, CompOut_F1, REGofMAX1DataOut_F1_46 ); 
OneRegister MUX1_F1_RO47(clk, write2_48, CompOut_F1, REGofMAX1DataOut_F1_47 ); 
OneRegister MUX1_F1_RO48(clk, write2_49, CompOut_F1, REGofMAX1DataOut_F1_48 ); 
OneRegister MUX1_F1_RO49(clk, write2_50, CompOut_F1, REGofMAX1DataOut_F1_49 ); 
OneRegister MUX1_F1_RO50(clk, write2_51, CompOut_F1, REGofMAX1DataOut_F1_50 ); 
OneRegister MUX1_F1_RO51(clk, write2_52, CompOut_F1, REGofMAX1DataOut_F1_51 ); 
OneRegister MUX1_F1_RO52(clk, write2_53, CompOut_F1, REGofMAX1DataOut_F1_52 ); 
OneRegister MUX1_F1_RO53(clk, write2_54, CompOut_F1, REGofMAX1DataOut_F1_53 ); 
OneRegister MUX1_F1_RO54(clk, write2_55, CompOut_F1, REGofMAX1DataOut_F1_54 ); 
OneRegister MUX1_F1_RO55(clk, write2_56, CompOut_F1, REGofMAX1DataOut_F1_55 ); 
OneRegister MUX1_F1_RO56(clk, write2_57, CompOut_F1, REGofMAX1DataOut_F1_56 ); 
OneRegister MUX1_F1_RO57(clk, write2_58, CompOut_F1, REGofMAX1DataOut_F1_57 ); 
OneRegister MUX1_F1_RO58(clk, write2_59, CompOut_F1, REGofMAX1DataOut_F1_58 ); 
OneRegister MUX1_F1_RO59(clk, write2_60, CompOut_F1, REGofMAX1DataOut_F1_59 ); 
OneRegister MUX1_F1_RO60(clk, write2_61, CompOut_F1, REGofMAX1DataOut_F1_60 ); 
OneRegister MUX1_F1_RO61(clk, write2_62, CompOut_F1, REGofMAX1DataOut_F1_61 ); 
OneRegister MUX1_F1_RO62(clk, write2_63, CompOut_F1, REGofMAX1DataOut_F1_62 ); 
OneRegister MUX1_F1_RO63(clk, write2_64, CompOut_F1, REGofMAX1DataOut_F1_63 ); 
OneRegister MUX1_F1_RO64(clk, write2_65, CompOut_F1, REGofMAX1DataOut_F1_64 ); 
OneRegister MUX1_F1_RO65(clk, write2_66, CompOut_F1, REGofMAX1DataOut_F1_65 ); 
OneRegister MUX1_F1_RO66(clk, write2_67, CompOut_F1, REGofMAX1DataOut_F1_66 ); 
OneRegister MUX1_F1_RO67(clk, write2_68, CompOut_F1, REGofMAX1DataOut_F1_67 ); 
OneRegister MUX1_F1_RO68(clk, write2_69, CompOut_F1, REGofMAX1DataOut_F1_68 ); 
OneRegister MUX1_F1_RO69(clk, write2_70, CompOut_F1, REGofMAX1DataOut_F1_69 ); 
OneRegister MUX1_F1_RO70(clk, write2_71, CompOut_F1, REGofMAX1DataOut_F1_70 ); 
OneRegister MUX1_F1_RO71(clk, write2_72, CompOut_F1, REGofMAX1DataOut_F1_71 ); 
OneRegister MUX1_F1_RO72(clk, write2_73, CompOut_F1, REGofMAX1DataOut_F1_72 ); 
OneRegister MUX1_F1_RO73(clk, write2_74, CompOut_F1, REGofMAX1DataOut_F1_73 ); 
OneRegister MUX1_F1_RO74(clk, write2_75, CompOut_F1, REGofMAX1DataOut_F1_74 ); 
OneRegister MUX1_F1_RO75(clk, write2_76, CompOut_F1, REGofMAX1DataOut_F1_75 ); 
OneRegister MUX1_F1_RO76(clk, write2_77, CompOut_F1, REGofMAX1DataOut_F1_76 ); 
OneRegister MUX1_F1_RO77(clk, write2_78, CompOut_F1, REGofMAX1DataOut_F1_77 ); 
OneRegister MUX1_F1_RO78(clk, write2_79, CompOut_F1, REGofMAX1DataOut_F1_78 ); 
OneRegister MUX1_F1_RO79(clk, write2_80, CompOut_F1, REGofMAX1DataOut_F1_79 ); 
OneRegister MUX1_F1_RO80(clk, write2_81, CompOut_F1, REGofMAX1DataOut_F1_80 ); 
OneRegister MUX1_F1_RO81(clk, write2_82, CompOut_F1, REGofMAX1DataOut_F1_81 ); 
OneRegister MUX1_F1_RO82(clk, write2_83, CompOut_F1, REGofMAX1DataOut_F1_82 ); 
OneRegister MUX1_F1_RO83(clk, write2_84, CompOut_F1, REGofMAX1DataOut_F1_83 ); 
OneRegister MUX1_F1_RO84(clk, write2_85, CompOut_F1, REGofMAX1DataOut_F1_84 ); 
OneRegister MUX1_F1_RO85(clk, write2_86, CompOut_F1, REGofMAX1DataOut_F1_85 ); 
OneRegister MUX1_F1_RO86(clk, write2_87, CompOut_F1, REGofMAX1DataOut_F1_86 ); 
OneRegister MUX1_F1_RO87(clk, write2_88, CompOut_F1, REGofMAX1DataOut_F1_87 ); 
OneRegister MUX1_F1_RO88(clk, write2_89, CompOut_F1, REGofMAX1DataOut_F1_88 ); 
OneRegister MUX1_F1_RO89(clk, write2_90, CompOut_F1, REGofMAX1DataOut_F1_89 ); 
OneRegister MUX1_F1_RO90(clk, write2_91, CompOut_F1, REGofMAX1DataOut_F1_90 ); 
OneRegister MUX1_F1_RO91(clk, write2_92, CompOut_F1, REGofMAX1DataOut_F1_91 ); 
OneRegister MUX1_F1_RO92(clk, write2_93, CompOut_F1, REGofMAX1DataOut_F1_92 ); 
OneRegister MUX1_F1_RO93(clk, write2_94, CompOut_F1, REGofMAX1DataOut_F1_93 ); 
OneRegister MUX1_F1_RO94(clk, write2_95, CompOut_F1, REGofMAX1DataOut_F1_94 ); 
OneRegister MUX1_F1_RO95(clk, write2_96, CompOut_F1, REGofMAX1DataOut_F1_95 ); 
OneRegister MUX1_F1_RO96(clk, write2_97, CompOut_F1, REGofMAX1DataOut_F1_96 ); 
OneRegister MUX1_F1_RO97(clk, write2_98, CompOut_F1, REGofMAX1DataOut_F1_97 ); 
OneRegister MUX1_F1_RO98(clk, write2_99, CompOut_F1, REGofMAX1DataOut_F1_98 ); 
OneRegister MUX1_F1_RO99(clk, write2_100, CompOut_F1, REGofMAX1DataOut_F1_99 ); 
OneRegister MUX1_F1_RO100(clk, write2_101, CompOut_F1, REGofMAX1DataOut_F1_100 ); 
OneRegister MUX1_F1_RO101(clk, write2_102, CompOut_F1, REGofMAX1DataOut_F1_101 ); 
OneRegister MUX1_F1_RO102(clk, write2_103, CompOut_F1, REGofMAX1DataOut_F1_102 ); 
OneRegister MUX1_F1_RO103(clk, write2_104, CompOut_F1, REGofMAX1DataOut_F1_103 ); 
OneRegister MUX1_F1_RO104(clk, write2_105, CompOut_F1, REGofMAX1DataOut_F1_104 ); 
OneRegister MUX1_F1_RO105(clk, write2_106, CompOut_F1, REGofMAX1DataOut_F1_105 ); 
OneRegister MUX1_F1_RO106(clk, write2_107, CompOut_F1, REGofMAX1DataOut_F1_106 ); 
OneRegister MUX1_F1_RO107(clk, write2_108, CompOut_F1, REGofMAX1DataOut_F1_107 ); 
OneRegister MUX1_F1_RO108(clk, write2_109, CompOut_F1, REGofMAX1DataOut_F1_108 ); 
OneRegister MUX1_F1_RO109(clk, write2_110, CompOut_F1, REGofMAX1DataOut_F1_109 ); 
OneRegister MUX1_F1_RO110(clk, write2_111, CompOut_F1, REGofMAX1DataOut_F1_110 ); 
OneRegister MUX1_F1_RO111(clk, write2_112, CompOut_F1, REGofMAX1DataOut_F1_111 ); 
OneRegister MUX1_F1_RO112(clk, write2_113, CompOut_F1, REGofMAX1DataOut_F1_112 ); 
OneRegister MUX1_F1_RO113(clk, write2_114, CompOut_F1, REGofMAX1DataOut_F1_113 ); 
OneRegister MUX1_F1_RO114(clk, write2_115, CompOut_F1, REGofMAX1DataOut_F1_114 ); 
OneRegister MUX1_F1_RO115(clk, write2_116, CompOut_F1, REGofMAX1DataOut_F1_115 ); 
OneRegister MUX1_F1_RO116(clk, write2_117, CompOut_F1, REGofMAX1DataOut_F1_116 ); 
OneRegister MUX1_F1_RO117(clk, write2_118, CompOut_F1, REGofMAX1DataOut_F1_117 ); 
OneRegister MUX1_F1_RO118(clk, write2_119, CompOut_F1, REGofMAX1DataOut_F1_118 ); 
OneRegister MUX1_F1_RO119(clk, write2_120, CompOut_F1, REGofMAX1DataOut_F1_119 ); 
OneRegister MUX1_F1_RO120(clk, write2_121, CompOut_F1, REGofMAX1DataOut_F1_120 ); 
OneRegister MUX1_F1_RO121(clk, write2_122, CompOut_F1, REGofMAX1DataOut_F1_121 ); 
OneRegister MUX1_F1_RO122(clk, write2_123, CompOut_F1, REGofMAX1DataOut_F1_122 ); 
OneRegister MUX1_F1_RO123(clk, write2_124, CompOut_F1, REGofMAX1DataOut_F1_123 ); 
OneRegister MUX1_F1_RO124(clk, write2_125, CompOut_F1, REGofMAX1DataOut_F1_124 ); 
OneRegister MUX1_F1_RO125(clk, write2_126, CompOut_F1, REGofMAX1DataOut_F1_125 ); 
OneRegister MUX1_F1_RO126(clk, write2_127, CompOut_F1, REGofMAX1DataOut_F1_126 ); 
OneRegister MUX1_F1_RO127(clk, write2_128, CompOut_F1, REGofMAX1DataOut_F1_127 ); 
OneRegister MUX1_F1_RO128(clk, write2_129, CompOut_F1, REGofMAX1DataOut_F1_128 ); 
OneRegister MUX1_F1_RO129(clk, write2_130, CompOut_F1, REGofMAX1DataOut_F1_129 ); 
OneRegister MUX1_F1_RO130(clk, write2_131, CompOut_F1, REGofMAX1DataOut_F1_130 ); 
OneRegister MUX1_F1_RO131(clk, write2_132, CompOut_F1, REGofMAX1DataOut_F1_131 ); 
OneRegister MUX1_F1_RO132(clk, write2_133, CompOut_F1, REGofMAX1DataOut_F1_132 ); 
OneRegister MUX1_F1_RO133(clk, write2_134, CompOut_F1, REGofMAX1DataOut_F1_133 ); 
OneRegister MUX1_F1_RO134(clk, write2_135, CompOut_F1, REGofMAX1DataOut_F1_134 ); 
OneRegister MUX1_F1_RO135(clk, write2_136, CompOut_F1, REGofMAX1DataOut_F1_135 ); 
OneRegister MUX1_F1_RO136(clk, write2_137, CompOut_F1, REGofMAX1DataOut_F1_136 ); 
OneRegister MUX1_F1_RO137(clk, write2_138, CompOut_F1, REGofMAX1DataOut_F1_137 ); 
OneRegister MUX1_F1_RO138(clk, write2_139, CompOut_F1, REGofMAX1DataOut_F1_138 ); 
OneRegister MUX1_F1_RO139(clk, write2_140, CompOut_F1, REGofMAX1DataOut_F1_139 ); 
OneRegister MUX1_F1_RO140(clk, write2_141, CompOut_F1, REGofMAX1DataOut_F1_140 ); 
OneRegister MUX1_F1_RO141(clk, write2_142, CompOut_F1, REGofMAX1DataOut_F1_141 ); 
OneRegister MUX1_F1_RO142(clk, write2_143, CompOut_F1, REGofMAX1DataOut_F1_142 ); 
OneRegister MUX1_F1_RO143(clk, write2_144, CompOut_F1, REGofMAX1DataOut_F1_143 ); 


///




OneRegister MUX1_F2_RO0(clk, write2_1, CompOut_F2, REGofMAX1DataOut_F2_0 ); 
OneRegister MUX1_F2_RO1(clk, write2_2, CompOut_F2, REGofMAX1DataOut_F2_1 ); 
OneRegister MUX1_F2_RO2(clk, write2_3, CompOut_F2, REGofMAX1DataOut_F2_2 ); 
OneRegister MUX1_F2_RO3(clk, write2_4, CompOut_F2, REGofMAX1DataOut_F2_3 ); 
OneRegister MUX1_F2_RO4(clk, write2_5, CompOut_F2, REGofMAX1DataOut_F2_4 ); 
OneRegister MUX1_F2_RO5(clk, write2_6, CompOut_F2, REGofMAX1DataOut_F2_5 ); 
OneRegister MUX1_F2_RO6(clk, write2_7, CompOut_F2, REGofMAX1DataOut_F2_6 ); 
OneRegister MUX1_F2_RO7(clk, write2_8, CompOut_F2, REGofMAX1DataOut_F2_7 ); 
OneRegister MUX1_F2_RO8(clk, write2_9, CompOut_F2, REGofMAX1DataOut_F2_8 ); 
OneRegister MUX1_F2_RO9(clk, write2_10, CompOut_F2, REGofMAX1DataOut_F2_9 ); 
OneRegister MUX1_F2_RO10(clk, write2_11, CompOut_F2, REGofMAX1DataOut_F2_10 ); 
OneRegister MUX1_F2_RO11(clk, write2_12, CompOut_F2, REGofMAX1DataOut_F2_11 ); 
OneRegister MUX1_F2_RO12(clk, write2_13, CompOut_F2, REGofMAX1DataOut_F2_12 ); 
OneRegister MUX1_F2_RO13(clk, write2_14, CompOut_F2, REGofMAX1DataOut_F2_13 ); 
OneRegister MUX1_F2_RO14(clk, write2_15, CompOut_F2, REGofMAX1DataOut_F2_14 ); 
OneRegister MUX1_F2_RO15(clk, write2_16, CompOut_F2, REGofMAX1DataOut_F2_15 ); 
OneRegister MUX1_F2_RO16(clk, write2_17, CompOut_F2, REGofMAX1DataOut_F2_16 ); 
OneRegister MUX1_F2_RO17(clk, write2_18, CompOut_F2, REGofMAX1DataOut_F2_17 ); 
OneRegister MUX1_F2_RO18(clk, write2_19, CompOut_F2, REGofMAX1DataOut_F2_18 ); 
OneRegister MUX1_F2_RO19(clk, write2_20, CompOut_F2, REGofMAX1DataOut_F2_19 ); 
OneRegister MUX1_F2_RO20(clk, write2_21, CompOut_F2, REGofMAX1DataOut_F2_20 ); 
OneRegister MUX1_F2_RO21(clk, write2_22, CompOut_F2, REGofMAX1DataOut_F2_21 ); 
OneRegister MUX1_F2_RO22(clk, write2_23, CompOut_F2, REGofMAX1DataOut_F2_22 ); 
OneRegister MUX1_F2_RO23(clk, write2_24, CompOut_F2, REGofMAX1DataOut_F2_23 ); 
OneRegister MUX1_F2_RO24(clk, write2_25, CompOut_F2, REGofMAX1DataOut_F2_24 ); 
OneRegister MUX1_F2_RO25(clk, write2_26, CompOut_F2, REGofMAX1DataOut_F2_25 ); 
OneRegister MUX1_F2_RO26(clk, write2_27, CompOut_F2, REGofMAX1DataOut_F2_26 ); 
OneRegister MUX1_F2_RO27(clk, write2_28, CompOut_F2, REGofMAX1DataOut_F2_27 ); 
OneRegister MUX1_F2_RO28(clk, write2_29, CompOut_F2, REGofMAX1DataOut_F2_28 ); 
OneRegister MUX1_F2_RO29(clk, write2_30, CompOut_F2, REGofMAX1DataOut_F2_29 ); 
OneRegister MUX1_F2_RO30(clk, write2_31, CompOut_F2, REGofMAX1DataOut_F2_30 ); 
OneRegister MUX1_F2_RO31(clk, write2_32, CompOut_F2, REGofMAX1DataOut_F2_31 ); 
OneRegister MUX1_F2_RO32(clk, write2_33, CompOut_F2, REGofMAX1DataOut_F2_32 ); 
OneRegister MUX1_F2_RO33(clk, write2_34, CompOut_F2, REGofMAX1DataOut_F2_33 ); 
OneRegister MUX1_F2_RO34(clk, write2_35, CompOut_F2, REGofMAX1DataOut_F2_34 ); 
OneRegister MUX1_F2_RO35(clk, write2_36, CompOut_F2, REGofMAX1DataOut_F2_35 ); 
OneRegister MUX1_F2_RO36(clk, write2_37, CompOut_F2, REGofMAX1DataOut_F2_36 ); 
OneRegister MUX1_F2_RO37(clk, write2_38, CompOut_F2, REGofMAX1DataOut_F2_37 ); 
OneRegister MUX1_F2_RO38(clk, write2_39, CompOut_F2, REGofMAX1DataOut_F2_38 ); 
OneRegister MUX1_F2_RO39(clk, write2_40, CompOut_F2, REGofMAX1DataOut_F2_39 ); 
OneRegister MUX1_F2_RO40(clk, write2_41, CompOut_F2, REGofMAX1DataOut_F2_40 ); 
OneRegister MUX1_F2_RO41(clk, write2_42, CompOut_F2, REGofMAX1DataOut_F2_41 ); 
OneRegister MUX1_F2_RO42(clk, write2_43, CompOut_F2, REGofMAX1DataOut_F2_42 ); 
OneRegister MUX1_F2_RO43(clk, write2_44, CompOut_F2, REGofMAX1DataOut_F2_43 ); 
OneRegister MUX1_F2_RO44(clk, write2_45, CompOut_F2, REGofMAX1DataOut_F2_44 ); 
OneRegister MUX1_F2_RO45(clk, write2_46, CompOut_F2, REGofMAX1DataOut_F2_45 ); 
OneRegister MUX1_F2_RO46(clk, write2_47, CompOut_F2, REGofMAX1DataOut_F2_46 ); 
OneRegister MUX1_F2_RO47(clk, write2_48, CompOut_F2, REGofMAX1DataOut_F2_47 ); 
OneRegister MUX1_F2_RO48(clk, write2_49, CompOut_F2, REGofMAX1DataOut_F2_48 ); 
OneRegister MUX1_F2_RO49(clk, write2_50, CompOut_F2, REGofMAX1DataOut_F2_49 ); 
OneRegister MUX1_F2_RO50(clk, write2_51, CompOut_F2, REGofMAX1DataOut_F2_50 ); 
OneRegister MUX1_F2_RO51(clk, write2_52, CompOut_F2, REGofMAX1DataOut_F2_51 ); 
OneRegister MUX1_F2_RO52(clk, write2_53, CompOut_F2, REGofMAX1DataOut_F2_52 ); 
OneRegister MUX1_F2_RO53(clk, write2_54, CompOut_F2, REGofMAX1DataOut_F2_53 ); 
OneRegister MUX1_F2_RO54(clk, write2_55, CompOut_F2, REGofMAX1DataOut_F2_54 ); 
OneRegister MUX1_F2_RO55(clk, write2_56, CompOut_F2, REGofMAX1DataOut_F2_55 ); 
OneRegister MUX1_F2_RO56(clk, write2_57, CompOut_F2, REGofMAX1DataOut_F2_56 ); 
OneRegister MUX1_F2_RO57(clk, write2_58, CompOut_F2, REGofMAX1DataOut_F2_57 ); 
OneRegister MUX1_F2_RO58(clk, write2_59, CompOut_F2, REGofMAX1DataOut_F2_58 ); 
OneRegister MUX1_F2_RO59(clk, write2_60, CompOut_F2, REGofMAX1DataOut_F2_59 ); 
OneRegister MUX1_F2_RO60(clk, write2_61, CompOut_F2, REGofMAX1DataOut_F2_60 ); 
OneRegister MUX1_F2_RO61(clk, write2_62, CompOut_F2, REGofMAX1DataOut_F2_61 ); 
OneRegister MUX1_F2_RO62(clk, write2_63, CompOut_F2, REGofMAX1DataOut_F2_62 ); 
OneRegister MUX1_F2_RO63(clk, write2_64, CompOut_F2, REGofMAX1DataOut_F2_63 ); 
OneRegister MUX1_F2_RO64(clk, write2_65, CompOut_F2, REGofMAX1DataOut_F2_64 ); 
OneRegister MUX1_F2_RO65(clk, write2_66, CompOut_F2, REGofMAX1DataOut_F2_65 ); 
OneRegister MUX1_F2_RO66(clk, write2_67, CompOut_F2, REGofMAX1DataOut_F2_66 ); 
OneRegister MUX1_F2_RO67(clk, write2_68, CompOut_F2, REGofMAX1DataOut_F2_67 ); 
OneRegister MUX1_F2_RO68(clk, write2_69, CompOut_F2, REGofMAX1DataOut_F2_68 ); 
OneRegister MUX1_F2_RO69(clk, write2_70, CompOut_F2, REGofMAX1DataOut_F2_69 ); 
OneRegister MUX1_F2_RO70(clk, write2_71, CompOut_F2, REGofMAX1DataOut_F2_70 ); 
OneRegister MUX1_F2_RO71(clk, write2_72, CompOut_F2, REGofMAX1DataOut_F2_71 ); 
OneRegister MUX1_F2_RO72(clk, write2_73, CompOut_F2, REGofMAX1DataOut_F2_72 ); 
OneRegister MUX1_F2_RO73(clk, write2_74, CompOut_F2, REGofMAX1DataOut_F2_73 ); 
OneRegister MUX1_F2_RO74(clk, write2_75, CompOut_F2, REGofMAX1DataOut_F2_74 ); 
OneRegister MUX1_F2_RO75(clk, write2_76, CompOut_F2, REGofMAX1DataOut_F2_75 ); 
OneRegister MUX1_F2_RO76(clk, write2_77, CompOut_F2, REGofMAX1DataOut_F2_76 ); 
OneRegister MUX1_F2_RO77(clk, write2_78, CompOut_F2, REGofMAX1DataOut_F2_77 ); 
OneRegister MUX1_F2_RO78(clk, write2_79, CompOut_F2, REGofMAX1DataOut_F2_78 ); 
OneRegister MUX1_F2_RO79(clk, write2_80, CompOut_F2, REGofMAX1DataOut_F2_79 ); 
OneRegister MUX1_F2_RO80(clk, write2_81, CompOut_F2, REGofMAX1DataOut_F2_80 ); 
OneRegister MUX1_F2_RO81(clk, write2_82, CompOut_F2, REGofMAX1DataOut_F2_81 ); 
OneRegister MUX1_F2_RO82(clk, write2_83, CompOut_F2, REGofMAX1DataOut_F2_82 ); 
OneRegister MUX1_F2_RO83(clk, write2_84, CompOut_F2, REGofMAX1DataOut_F2_83 ); 
OneRegister MUX1_F2_RO84(clk, write2_85, CompOut_F2, REGofMAX1DataOut_F2_84 ); 
OneRegister MUX1_F2_RO85(clk, write2_86, CompOut_F2, REGofMAX1DataOut_F2_85 ); 
OneRegister MUX1_F2_RO86(clk, write2_87, CompOut_F2, REGofMAX1DataOut_F2_86 ); 
OneRegister MUX1_F2_RO87(clk, write2_88, CompOut_F2, REGofMAX1DataOut_F2_87 ); 
OneRegister MUX1_F2_RO88(clk, write2_89, CompOut_F2, REGofMAX1DataOut_F2_88 ); 
OneRegister MUX1_F2_RO89(clk, write2_90, CompOut_F2, REGofMAX1DataOut_F2_89 ); 
OneRegister MUX1_F2_RO90(clk, write2_91, CompOut_F2, REGofMAX1DataOut_F2_90 ); 
OneRegister MUX1_F2_RO91(clk, write2_92, CompOut_F2, REGofMAX1DataOut_F2_91 ); 
OneRegister MUX1_F2_RO92(clk, write2_93, CompOut_F2, REGofMAX1DataOut_F2_92 ); 
OneRegister MUX1_F2_RO93(clk, write2_94, CompOut_F2, REGofMAX1DataOut_F2_93 ); 
OneRegister MUX1_F2_RO94(clk, write2_95, CompOut_F2, REGofMAX1DataOut_F2_94 ); 
OneRegister MUX1_F2_RO95(clk, write2_96, CompOut_F2, REGofMAX1DataOut_F2_95 ); 
OneRegister MUX1_F2_RO96(clk, write2_97, CompOut_F2, REGofMAX1DataOut_F2_96 ); 
OneRegister MUX1_F2_RO97(clk, write2_98, CompOut_F2, REGofMAX1DataOut_F2_97 ); 
OneRegister MUX1_F2_RO98(clk, write2_99, CompOut_F2, REGofMAX1DataOut_F2_98 ); 
OneRegister MUX1_F2_RO99(clk, write2_100, CompOut_F2, REGofMAX1DataOut_F2_99 ); 
OneRegister MUX1_F2_RO100(clk, write2_101, CompOut_F2, REGofMAX1DataOut_F2_100 ); 
OneRegister MUX1_F2_RO101(clk, write2_102, CompOut_F2, REGofMAX1DataOut_F2_101 ); 
OneRegister MUX1_F2_RO102(clk, write2_103, CompOut_F2, REGofMAX1DataOut_F2_102 ); 
OneRegister MUX1_F2_RO103(clk, write2_104, CompOut_F2, REGofMAX1DataOut_F2_103 ); 
OneRegister MUX1_F2_RO104(clk, write2_105, CompOut_F2, REGofMAX1DataOut_F2_104 ); 
OneRegister MUX1_F2_RO105(clk, write2_106, CompOut_F2, REGofMAX1DataOut_F2_105 ); 
OneRegister MUX1_F2_RO106(clk, write2_107, CompOut_F2, REGofMAX1DataOut_F2_106 ); 
OneRegister MUX1_F2_RO107(clk, write2_108, CompOut_F2, REGofMAX1DataOut_F2_107 ); 
OneRegister MUX1_F2_RO108(clk, write2_109, CompOut_F2, REGofMAX1DataOut_F2_108 ); 
OneRegister MUX1_F2_RO109(clk, write2_110, CompOut_F2, REGofMAX1DataOut_F2_109 ); 
OneRegister MUX1_F2_RO110(clk, write2_111, CompOut_F2, REGofMAX1DataOut_F2_110 ); 
OneRegister MUX1_F2_RO111(clk, write2_112, CompOut_F2, REGofMAX1DataOut_F2_111 ); 
OneRegister MUX1_F2_RO112(clk, write2_113, CompOut_F2, REGofMAX1DataOut_F2_112 ); 
OneRegister MUX1_F2_RO113(clk, write2_114, CompOut_F2, REGofMAX1DataOut_F2_113 ); 
OneRegister MUX1_F2_RO114(clk, write2_115, CompOut_F2, REGofMAX1DataOut_F2_114 ); 
OneRegister MUX1_F2_RO115(clk, write2_116, CompOut_F2, REGofMAX1DataOut_F2_115 ); 
OneRegister MUX1_F2_RO116(clk, write2_117, CompOut_F2, REGofMAX1DataOut_F2_116 ); 
OneRegister MUX1_F2_RO117(clk, write2_118, CompOut_F2, REGofMAX1DataOut_F2_117 ); 
OneRegister MUX1_F2_RO118(clk, write2_119, CompOut_F2, REGofMAX1DataOut_F2_118 ); 
OneRegister MUX1_F2_RO119(clk, write2_120, CompOut_F2, REGofMAX1DataOut_F2_119 ); 
OneRegister MUX1_F2_RO120(clk, write2_121, CompOut_F2, REGofMAX1DataOut_F2_120 ); 
OneRegister MUX1_F2_RO121(clk, write2_122, CompOut_F2, REGofMAX1DataOut_F2_121 ); 
OneRegister MUX1_F2_RO122(clk, write2_123, CompOut_F2, REGofMAX1DataOut_F2_122 ); 
OneRegister MUX1_F2_RO123(clk, write2_124, CompOut_F2, REGofMAX1DataOut_F2_123 ); 
OneRegister MUX1_F2_RO124(clk, write2_125, CompOut_F2, REGofMAX1DataOut_F2_124 ); 
OneRegister MUX1_F2_RO125(clk, write2_126, CompOut_F2, REGofMAX1DataOut_F2_125 ); 
OneRegister MUX1_F2_RO126(clk, write2_127, CompOut_F2, REGofMAX1DataOut_F2_126 ); 
OneRegister MUX1_F2_RO127(clk, write2_128, CompOut_F2, REGofMAX1DataOut_F2_127 ); 
OneRegister MUX1_F2_RO128(clk, write2_129, CompOut_F2, REGofMAX1DataOut_F2_128 ); 
OneRegister MUX1_F2_RO129(clk, write2_130, CompOut_F2, REGofMAX1DataOut_F2_129 ); 
OneRegister MUX1_F2_RO130(clk, write2_131, CompOut_F2, REGofMAX1DataOut_F2_130 ); 
OneRegister MUX1_F2_RO131(clk, write2_132, CompOut_F2, REGofMAX1DataOut_F2_131 ); 
OneRegister MUX1_F2_RO132(clk, write2_133, CompOut_F2, REGofMAX1DataOut_F2_132 ); 
OneRegister MUX1_F2_RO133(clk, write2_134, CompOut_F2, REGofMAX1DataOut_F2_133 ); 
OneRegister MUX1_F2_RO134(clk, write2_135, CompOut_F2, REGofMAX1DataOut_F2_134 ); 
OneRegister MUX1_F2_RO135(clk, write2_136, CompOut_F2, REGofMAX1DataOut_F2_135 ); 
OneRegister MUX1_F2_RO136(clk, write2_137, CompOut_F2, REGofMAX1DataOut_F2_136 ); 
OneRegister MUX1_F2_RO137(clk, write2_138, CompOut_F2, REGofMAX1DataOut_F2_137 ); 
OneRegister MUX1_F2_RO138(clk, write2_139, CompOut_F2, REGofMAX1DataOut_F2_138 ); 
OneRegister MUX1_F2_RO139(clk, write2_140, CompOut_F2, REGofMAX1DataOut_F2_139 ); 
OneRegister MUX1_F2_RO140(clk, write2_141, CompOut_F2, REGofMAX1DataOut_F2_140 ); 
OneRegister MUX1_F2_RO141(clk, write2_142, CompOut_F2, REGofMAX1DataOut_F2_141 ); 
OneRegister MUX1_F2_RO142(clk, write2_143, CompOut_F2, REGofMAX1DataOut_F2_142 ); 
OneRegister MUX1_F2_RO143(clk, write2_144, CompOut_F2, REGofMAX1DataOut_F2_143 ); 

///



OneRegister MUX1_F3_RO0(clk, write2_1, CompOut_F3, REGofMAX1DataOut_F3_0 ); 
OneRegister MUX1_F3_RO1(clk, write2_2, CompOut_F3, REGofMAX1DataOut_F3_1 ); 
OneRegister MUX1_F3_RO2(clk, write2_3, CompOut_F3, REGofMAX1DataOut_F3_2 ); 
OneRegister MUX1_F3_RO3(clk, write2_4, CompOut_F3, REGofMAX1DataOut_F3_3 ); 
OneRegister MUX1_F3_RO4(clk, write2_5, CompOut_F3, REGofMAX1DataOut_F3_4 ); 
OneRegister MUX1_F3_RO5(clk, write2_6, CompOut_F3, REGofMAX1DataOut_F3_5 ); 
OneRegister MUX1_F3_RO6(clk, write2_7, CompOut_F3, REGofMAX1DataOut_F3_6 ); 
OneRegister MUX1_F3_RO7(clk, write2_8, CompOut_F3, REGofMAX1DataOut_F3_7 ); 
OneRegister MUX1_F3_RO8(clk, write2_9, CompOut_F3, REGofMAX1DataOut_F3_8 ); 
OneRegister MUX1_F3_RO9(clk, write2_10, CompOut_F3, REGofMAX1DataOut_F3_9 ); 
OneRegister MUX1_F3_RO10(clk, write2_11, CompOut_F3, REGofMAX1DataOut_F3_10 ); 
OneRegister MUX1_F3_RO11(clk, write2_12, CompOut_F3, REGofMAX1DataOut_F3_11 ); 
OneRegister MUX1_F3_RO12(clk, write2_13, CompOut_F3, REGofMAX1DataOut_F3_12 ); 
OneRegister MUX1_F3_RO13(clk, write2_14, CompOut_F3, REGofMAX1DataOut_F3_13 ); 
OneRegister MUX1_F3_RO14(clk, write2_15, CompOut_F3, REGofMAX1DataOut_F3_14 ); 
OneRegister MUX1_F3_RO15(clk, write2_16, CompOut_F3, REGofMAX1DataOut_F3_15 ); 
OneRegister MUX1_F3_RO16(clk, write2_17, CompOut_F3, REGofMAX1DataOut_F3_16 ); 
OneRegister MUX1_F3_RO17(clk, write2_18, CompOut_F3, REGofMAX1DataOut_F3_17 ); 
OneRegister MUX1_F3_RO18(clk, write2_19, CompOut_F3, REGofMAX1DataOut_F3_18 ); 
OneRegister MUX1_F3_RO19(clk, write2_20, CompOut_F3, REGofMAX1DataOut_F3_19 ); 
OneRegister MUX1_F3_RO20(clk, write2_21, CompOut_F3, REGofMAX1DataOut_F3_20 ); 
OneRegister MUX1_F3_RO21(clk, write2_22, CompOut_F3, REGofMAX1DataOut_F3_21 ); 
OneRegister MUX1_F3_RO22(clk, write2_23, CompOut_F3, REGofMAX1DataOut_F3_22 ); 
OneRegister MUX1_F3_RO23(clk, write2_24, CompOut_F3, REGofMAX1DataOut_F3_23 ); 
OneRegister MUX1_F3_RO24(clk, write2_25, CompOut_F3, REGofMAX1DataOut_F3_24 ); 
OneRegister MUX1_F3_RO25(clk, write2_26, CompOut_F3, REGofMAX1DataOut_F3_25 ); 
OneRegister MUX1_F3_RO26(clk, write2_27, CompOut_F3, REGofMAX1DataOut_F3_26 ); 
OneRegister MUX1_F3_RO27(clk, write2_28, CompOut_F3, REGofMAX1DataOut_F3_27 ); 
OneRegister MUX1_F3_RO28(clk, write2_29, CompOut_F3, REGofMAX1DataOut_F3_28 ); 
OneRegister MUX1_F3_RO29(clk, write2_30, CompOut_F3, REGofMAX1DataOut_F3_29 ); 
OneRegister MUX1_F3_RO30(clk, write2_31, CompOut_F3, REGofMAX1DataOut_F3_30 ); 
OneRegister MUX1_F3_RO31(clk, write2_32, CompOut_F3, REGofMAX1DataOut_F3_31 ); 
OneRegister MUX1_F3_RO32(clk, write2_33, CompOut_F3, REGofMAX1DataOut_F3_32 ); 
OneRegister MUX1_F3_RO33(clk, write2_34, CompOut_F3, REGofMAX1DataOut_F3_33 ); 
OneRegister MUX1_F3_RO34(clk, write2_35, CompOut_F3, REGofMAX1DataOut_F3_34 ); 
OneRegister MUX1_F3_RO35(clk, write2_36, CompOut_F3, REGofMAX1DataOut_F3_35 ); 
OneRegister MUX1_F3_RO36(clk, write2_37, CompOut_F3, REGofMAX1DataOut_F3_36 ); 
OneRegister MUX1_F3_RO37(clk, write2_38, CompOut_F3, REGofMAX1DataOut_F3_37 ); 
OneRegister MUX1_F3_RO38(clk, write2_39, CompOut_F3, REGofMAX1DataOut_F3_38 ); 
OneRegister MUX1_F3_RO39(clk, write2_40, CompOut_F3, REGofMAX1DataOut_F3_39 ); 
OneRegister MUX1_F3_RO40(clk, write2_41, CompOut_F3, REGofMAX1DataOut_F3_40 ); 
OneRegister MUX1_F3_RO41(clk, write2_42, CompOut_F3, REGofMAX1DataOut_F3_41 ); 
OneRegister MUX1_F3_RO42(clk, write2_43, CompOut_F3, REGofMAX1DataOut_F3_42 ); 
OneRegister MUX1_F3_RO43(clk, write2_44, CompOut_F3, REGofMAX1DataOut_F3_43 ); 
OneRegister MUX1_F3_RO44(clk, write2_45, CompOut_F3, REGofMAX1DataOut_F3_44 ); 
OneRegister MUX1_F3_RO45(clk, write2_46, CompOut_F3, REGofMAX1DataOut_F3_45 ); 
OneRegister MUX1_F3_RO46(clk, write2_47, CompOut_F3, REGofMAX1DataOut_F3_46 ); 
OneRegister MUX1_F3_RO47(clk, write2_48, CompOut_F3, REGofMAX1DataOut_F3_47 ); 
OneRegister MUX1_F3_RO48(clk, write2_49, CompOut_F3, REGofMAX1DataOut_F3_48 ); 
OneRegister MUX1_F3_RO49(clk, write2_50, CompOut_F3, REGofMAX1DataOut_F3_49 ); 
OneRegister MUX1_F3_RO50(clk, write2_51, CompOut_F3, REGofMAX1DataOut_F3_50 ); 
OneRegister MUX1_F3_RO51(clk, write2_52, CompOut_F3, REGofMAX1DataOut_F3_51 ); 
OneRegister MUX1_F3_RO52(clk, write2_53, CompOut_F3, REGofMAX1DataOut_F3_52 ); 
OneRegister MUX1_F3_RO53(clk, write2_54, CompOut_F3, REGofMAX1DataOut_F3_53 ); 
OneRegister MUX1_F3_RO54(clk, write2_55, CompOut_F3, REGofMAX1DataOut_F3_54 ); 
OneRegister MUX1_F3_RO55(clk, write2_56, CompOut_F3, REGofMAX1DataOut_F3_55 ); 
OneRegister MUX1_F3_RO56(clk, write2_57, CompOut_F3, REGofMAX1DataOut_F3_56 ); 
OneRegister MUX1_F3_RO57(clk, write2_58, CompOut_F3, REGofMAX1DataOut_F3_57 ); 
OneRegister MUX1_F3_RO58(clk, write2_59, CompOut_F3, REGofMAX1DataOut_F3_58 ); 
OneRegister MUX1_F3_RO59(clk, write2_60, CompOut_F3, REGofMAX1DataOut_F3_59 ); 
OneRegister MUX1_F3_RO60(clk, write2_61, CompOut_F3, REGofMAX1DataOut_F3_60 ); 
OneRegister MUX1_F3_RO61(clk, write2_62, CompOut_F3, REGofMAX1DataOut_F3_61 ); 
OneRegister MUX1_F3_RO62(clk, write2_63, CompOut_F3, REGofMAX1DataOut_F3_62 ); 
OneRegister MUX1_F3_RO63(clk, write2_64, CompOut_F3, REGofMAX1DataOut_F3_63 ); 
OneRegister MUX1_F3_RO64(clk, write2_65, CompOut_F3, REGofMAX1DataOut_F3_64 ); 
OneRegister MUX1_F3_RO65(clk, write2_66, CompOut_F3, REGofMAX1DataOut_F3_65 ); 
OneRegister MUX1_F3_RO66(clk, write2_67, CompOut_F3, REGofMAX1DataOut_F3_66 ); 
OneRegister MUX1_F3_RO67(clk, write2_68, CompOut_F3, REGofMAX1DataOut_F3_67 ); 
OneRegister MUX1_F3_RO68(clk, write2_69, CompOut_F3, REGofMAX1DataOut_F3_68 ); 
OneRegister MUX1_F3_RO69(clk, write2_70, CompOut_F3, REGofMAX1DataOut_F3_69 ); 
OneRegister MUX1_F3_RO70(clk, write2_71, CompOut_F3, REGofMAX1DataOut_F3_70 ); 
OneRegister MUX1_F3_RO71(clk, write2_72, CompOut_F3, REGofMAX1DataOut_F3_71 ); 
OneRegister MUX1_F3_RO72(clk, write2_73, CompOut_F3, REGofMAX1DataOut_F3_72 ); 
OneRegister MUX1_F3_RO73(clk, write2_74, CompOut_F3, REGofMAX1DataOut_F3_73 ); 
OneRegister MUX1_F3_RO74(clk, write2_75, CompOut_F3, REGofMAX1DataOut_F3_74 ); 
OneRegister MUX1_F3_RO75(clk, write2_76, CompOut_F3, REGofMAX1DataOut_F3_75 ); 
OneRegister MUX1_F3_RO76(clk, write2_77, CompOut_F3, REGofMAX1DataOut_F3_76 ); 
OneRegister MUX1_F3_RO77(clk, write2_78, CompOut_F3, REGofMAX1DataOut_F3_77 ); 
OneRegister MUX1_F3_RO78(clk, write2_79, CompOut_F3, REGofMAX1DataOut_F3_78 ); 
OneRegister MUX1_F3_RO79(clk, write2_80, CompOut_F3, REGofMAX1DataOut_F3_79 ); 
OneRegister MUX1_F3_RO80(clk, write2_81, CompOut_F3, REGofMAX1DataOut_F3_80 ); 
OneRegister MUX1_F3_RO81(clk, write2_82, CompOut_F3, REGofMAX1DataOut_F3_81 ); 
OneRegister MUX1_F3_RO82(clk, write2_83, CompOut_F3, REGofMAX1DataOut_F3_82 ); 
OneRegister MUX1_F3_RO83(clk, write2_84, CompOut_F3, REGofMAX1DataOut_F3_83 ); 
OneRegister MUX1_F3_RO84(clk, write2_85, CompOut_F3, REGofMAX1DataOut_F3_84 ); 
OneRegister MUX1_F3_RO85(clk, write2_86, CompOut_F3, REGofMAX1DataOut_F3_85 ); 
OneRegister MUX1_F3_RO86(clk, write2_87, CompOut_F3, REGofMAX1DataOut_F3_86 ); 
OneRegister MUX1_F3_RO87(clk, write2_88, CompOut_F3, REGofMAX1DataOut_F3_87 ); 
OneRegister MUX1_F3_RO88(clk, write2_89, CompOut_F3, REGofMAX1DataOut_F3_88 ); 
OneRegister MUX1_F3_RO89(clk, write2_90, CompOut_F3, REGofMAX1DataOut_F3_89 ); 
OneRegister MUX1_F3_RO90(clk, write2_91, CompOut_F3, REGofMAX1DataOut_F3_90 ); 
OneRegister MUX1_F3_RO91(clk, write2_92, CompOut_F3, REGofMAX1DataOut_F3_91 ); 
OneRegister MUX1_F3_RO92(clk, write2_93, CompOut_F3, REGofMAX1DataOut_F3_92 ); 
OneRegister MUX1_F3_RO93(clk, write2_94, CompOut_F3, REGofMAX1DataOut_F3_93 ); 
OneRegister MUX1_F3_RO94(clk, write2_95, CompOut_F3, REGofMAX1DataOut_F3_94 ); 
OneRegister MUX1_F3_RO95(clk, write2_96, CompOut_F3, REGofMAX1DataOut_F3_95 ); 
OneRegister MUX1_F3_RO96(clk, write2_97, CompOut_F3, REGofMAX1DataOut_F3_96 ); 
OneRegister MUX1_F3_RO97(clk, write2_98, CompOut_F3, REGofMAX1DataOut_F3_97 ); 
OneRegister MUX1_F3_RO98(clk, write2_99, CompOut_F3, REGofMAX1DataOut_F3_98 ); 
OneRegister MUX1_F3_RO99(clk, write2_100, CompOut_F3, REGofMAX1DataOut_F3_99 ); 
OneRegister MUX1_F3_RO100(clk, write2_101, CompOut_F3, REGofMAX1DataOut_F3_100 ); 
OneRegister MUX1_F3_RO101(clk, write2_102, CompOut_F3, REGofMAX1DataOut_F3_101 ); 
OneRegister MUX1_F3_RO102(clk, write2_103, CompOut_F3, REGofMAX1DataOut_F3_102 ); 
OneRegister MUX1_F3_RO103(clk, write2_104, CompOut_F3, REGofMAX1DataOut_F3_103 ); 
OneRegister MUX1_F3_RO104(clk, write2_105, CompOut_F3, REGofMAX1DataOut_F3_104 ); 
OneRegister MUX1_F3_RO105(clk, write2_106, CompOut_F3, REGofMAX1DataOut_F3_105 ); 
OneRegister MUX1_F3_RO106(clk, write2_107, CompOut_F3, REGofMAX1DataOut_F3_106 ); 
OneRegister MUX1_F3_RO107(clk, write2_108, CompOut_F3, REGofMAX1DataOut_F3_107 ); 
OneRegister MUX1_F3_RO108(clk, write2_109, CompOut_F3, REGofMAX1DataOut_F3_108 ); 
OneRegister MUX1_F3_RO109(clk, write2_110, CompOut_F3, REGofMAX1DataOut_F3_109 ); 
OneRegister MUX1_F3_RO110(clk, write2_111, CompOut_F3, REGofMAX1DataOut_F3_110 ); 
OneRegister MUX1_F3_RO111(clk, write2_112, CompOut_F3, REGofMAX1DataOut_F3_111 ); 
OneRegister MUX1_F3_RO112(clk, write2_113, CompOut_F3, REGofMAX1DataOut_F3_112 ); 
OneRegister MUX1_F3_RO113(clk, write2_114, CompOut_F3, REGofMAX1DataOut_F3_113 ); 
OneRegister MUX1_F3_RO114(clk, write2_115, CompOut_F3, REGofMAX1DataOut_F3_114 ); 
OneRegister MUX1_F3_RO115(clk, write2_116, CompOut_F3, REGofMAX1DataOut_F3_115 ); 
OneRegister MUX1_F3_RO116(clk, write2_117, CompOut_F3, REGofMAX1DataOut_F3_116 ); 
OneRegister MUX1_F3_RO117(clk, write2_118, CompOut_F3, REGofMAX1DataOut_F3_117 ); 
OneRegister MUX1_F3_RO118(clk, write2_119, CompOut_F3, REGofMAX1DataOut_F3_118 ); 
OneRegister MUX1_F3_RO119(clk, write2_120, CompOut_F3, REGofMAX1DataOut_F3_119 ); 
OneRegister MUX1_F3_RO120(clk, write2_121, CompOut_F3, REGofMAX1DataOut_F3_120 ); 
OneRegister MUX1_F3_RO121(clk, write2_122, CompOut_F3, REGofMAX1DataOut_F3_121 ); 
OneRegister MUX1_F3_RO122(clk, write2_123, CompOut_F3, REGofMAX1DataOut_F3_122 ); 
OneRegister MUX1_F3_RO123(clk, write2_124, CompOut_F3, REGofMAX1DataOut_F3_123 ); 
OneRegister MUX1_F3_RO124(clk, write2_125, CompOut_F3, REGofMAX1DataOut_F3_124 ); 
OneRegister MUX1_F3_RO125(clk, write2_126, CompOut_F3, REGofMAX1DataOut_F3_125 ); 
OneRegister MUX1_F3_RO126(clk, write2_127, CompOut_F3, REGofMAX1DataOut_F3_126 ); 
OneRegister MUX1_F3_RO127(clk, write2_128, CompOut_F3, REGofMAX1DataOut_F3_127 ); 
OneRegister MUX1_F3_RO128(clk, write2_129, CompOut_F3, REGofMAX1DataOut_F3_128 ); 
OneRegister MUX1_F3_RO129(clk, write2_130, CompOut_F3, REGofMAX1DataOut_F3_129 ); 
OneRegister MUX1_F3_RO130(clk, write2_131, CompOut_F3, REGofMAX1DataOut_F3_130 ); 
OneRegister MUX1_F3_RO131(clk, write2_132, CompOut_F3, REGofMAX1DataOut_F3_131 ); 
OneRegister MUX1_F3_RO132(clk, write2_133, CompOut_F3, REGofMAX1DataOut_F3_132 ); 
OneRegister MUX1_F3_RO133(clk, write2_134, CompOut_F3, REGofMAX1DataOut_F3_133 ); 
OneRegister MUX1_F3_RO134(clk, write2_135, CompOut_F3, REGofMAX1DataOut_F3_134 ); 
OneRegister MUX1_F3_RO135(clk, write2_136, CompOut_F3, REGofMAX1DataOut_F3_135 ); 
OneRegister MUX1_F3_RO136(clk, write2_137, CompOut_F3, REGofMAX1DataOut_F3_136 ); 
OneRegister MUX1_F3_RO137(clk, write2_138, CompOut_F3, REGofMAX1DataOut_F3_137 ); 
OneRegister MUX1_F3_RO138(clk, write2_139, CompOut_F3, REGofMAX1DataOut_F3_138 ); 
OneRegister MUX1_F3_RO139(clk, write2_140, CompOut_F3, REGofMAX1DataOut_F3_139 ); 
OneRegister MUX1_F3_RO140(clk, write2_141, CompOut_F3, REGofMAX1DataOut_F3_140 ); 
OneRegister MUX1_F3_RO141(clk, write2_142, CompOut_F3, REGofMAX1DataOut_F3_141 ); 
OneRegister MUX1_F3_RO142(clk, write2_143, CompOut_F3, REGofMAX1DataOut_F3_142 ); 
OneRegister MUX1_F3_RO143(clk, write2_144, CompOut_F3, REGofMAX1DataOut_F3_143 ); 

//




OneRegister MUX1_F4_RO0(clk, write2_1, CompOut_F4, REGofMAX1DataOut_F4_0 ); 
OneRegister MUX1_F4_RO1(clk, write2_2, CompOut_F4, REGofMAX1DataOut_F4_1 ); 
OneRegister MUX1_F4_RO2(clk, write2_3, CompOut_F4, REGofMAX1DataOut_F4_2 ); 
OneRegister MUX1_F4_RO3(clk, write2_4, CompOut_F4, REGofMAX1DataOut_F4_3 ); 
OneRegister MUX1_F4_RO4(clk, write2_5, CompOut_F4, REGofMAX1DataOut_F4_4 ); 
OneRegister MUX1_F4_RO5(clk, write2_6, CompOut_F4, REGofMAX1DataOut_F4_5 ); 
OneRegister MUX1_F4_RO6(clk, write2_7, CompOut_F4, REGofMAX1DataOut_F4_6 ); 
OneRegister MUX1_F4_RO7(clk, write2_8, CompOut_F4, REGofMAX1DataOut_F4_7 ); 
OneRegister MUX1_F4_RO8(clk, write2_9, CompOut_F4, REGofMAX1DataOut_F4_8 ); 
OneRegister MUX1_F4_RO9(clk, write2_10, CompOut_F4, REGofMAX1DataOut_F4_9 ); 
OneRegister MUX1_F4_RO10(clk, write2_11, CompOut_F4, REGofMAX1DataOut_F4_10 ); 
OneRegister MUX1_F4_RO11(clk, write2_12, CompOut_F4, REGofMAX1DataOut_F4_11 ); 
OneRegister MUX1_F4_RO12(clk, write2_13, CompOut_F4, REGofMAX1DataOut_F4_12 ); 
OneRegister MUX1_F4_RO13(clk, write2_14, CompOut_F4, REGofMAX1DataOut_F4_13 ); 
OneRegister MUX1_F4_RO14(clk, write2_15, CompOut_F4, REGofMAX1DataOut_F4_14 ); 
OneRegister MUX1_F4_RO15(clk, write2_16, CompOut_F4, REGofMAX1DataOut_F4_15 ); 
OneRegister MUX1_F4_RO16(clk, write2_17, CompOut_F4, REGofMAX1DataOut_F4_16 ); 
OneRegister MUX1_F4_RO17(clk, write2_18, CompOut_F4, REGofMAX1DataOut_F4_17 ); 
OneRegister MUX1_F4_RO18(clk, write2_19, CompOut_F4, REGofMAX1DataOut_F4_18 ); 
OneRegister MUX1_F4_RO19(clk, write2_20, CompOut_F4, REGofMAX1DataOut_F4_19 ); 
OneRegister MUX1_F4_RO20(clk, write2_21, CompOut_F4, REGofMAX1DataOut_F4_20 ); 
OneRegister MUX1_F4_RO21(clk, write2_22, CompOut_F4, REGofMAX1DataOut_F4_21 ); 
OneRegister MUX1_F4_RO22(clk, write2_23, CompOut_F4, REGofMAX1DataOut_F4_22 ); 
OneRegister MUX1_F4_RO23(clk, write2_24, CompOut_F4, REGofMAX1DataOut_F4_23 ); 
OneRegister MUX1_F4_RO24(clk, write2_25, CompOut_F4, REGofMAX1DataOut_F4_24 ); 
OneRegister MUX1_F4_RO25(clk, write2_26, CompOut_F4, REGofMAX1DataOut_F4_25 ); 
OneRegister MUX1_F4_RO26(clk, write2_27, CompOut_F4, REGofMAX1DataOut_F4_26 ); 
OneRegister MUX1_F4_RO27(clk, write2_28, CompOut_F4, REGofMAX1DataOut_F4_27 ); 
OneRegister MUX1_F4_RO28(clk, write2_29, CompOut_F4, REGofMAX1DataOut_F4_28 ); 
OneRegister MUX1_F4_RO29(clk, write2_30, CompOut_F4, REGofMAX1DataOut_F4_29 ); 
OneRegister MUX1_F4_RO30(clk, write2_31, CompOut_F4, REGofMAX1DataOut_F4_30 ); 
OneRegister MUX1_F4_RO31(clk, write2_32, CompOut_F4, REGofMAX1DataOut_F4_31 ); 
OneRegister MUX1_F4_RO32(clk, write2_33, CompOut_F4, REGofMAX1DataOut_F4_32 ); 
OneRegister MUX1_F4_RO33(clk, write2_34, CompOut_F4, REGofMAX1DataOut_F4_33 ); 
OneRegister MUX1_F4_RO34(clk, write2_35, CompOut_F4, REGofMAX1DataOut_F4_34 ); 
OneRegister MUX1_F4_RO35(clk, write2_36, CompOut_F4, REGofMAX1DataOut_F4_35 ); 
OneRegister MUX1_F4_RO36(clk, write2_37, CompOut_F4, REGofMAX1DataOut_F4_36 ); 
OneRegister MUX1_F4_RO37(clk, write2_38, CompOut_F4, REGofMAX1DataOut_F4_37 ); 
OneRegister MUX1_F4_RO38(clk, write2_39, CompOut_F4, REGofMAX1DataOut_F4_38 ); 
OneRegister MUX1_F4_RO39(clk, write2_40, CompOut_F4, REGofMAX1DataOut_F4_39 ); 
OneRegister MUX1_F4_RO40(clk, write2_41, CompOut_F4, REGofMAX1DataOut_F4_40 ); 
OneRegister MUX1_F4_RO41(clk, write2_42, CompOut_F4, REGofMAX1DataOut_F4_41 ); 
OneRegister MUX1_F4_RO42(clk, write2_43, CompOut_F4, REGofMAX1DataOut_F4_42 ); 
OneRegister MUX1_F4_RO43(clk, write2_44, CompOut_F4, REGofMAX1DataOut_F4_43 ); 
OneRegister MUX1_F4_RO44(clk, write2_45, CompOut_F4, REGofMAX1DataOut_F4_44 ); 
OneRegister MUX1_F4_RO45(clk, write2_46, CompOut_F4, REGofMAX1DataOut_F4_45 ); 
OneRegister MUX1_F4_RO46(clk, write2_47, CompOut_F4, REGofMAX1DataOut_F4_46 ); 
OneRegister MUX1_F4_RO47(clk, write2_48, CompOut_F4, REGofMAX1DataOut_F4_47 ); 
OneRegister MUX1_F4_RO48(clk, write2_49, CompOut_F4, REGofMAX1DataOut_F4_48 ); 
OneRegister MUX1_F4_RO49(clk, write2_50, CompOut_F4, REGofMAX1DataOut_F4_49 ); 
OneRegister MUX1_F4_RO50(clk, write2_51, CompOut_F4, REGofMAX1DataOut_F4_50 ); 
OneRegister MUX1_F4_RO51(clk, write2_52, CompOut_F4, REGofMAX1DataOut_F4_51 ); 
OneRegister MUX1_F4_RO52(clk, write2_53, CompOut_F4, REGofMAX1DataOut_F4_52 ); 
OneRegister MUX1_F4_RO53(clk, write2_54, CompOut_F4, REGofMAX1DataOut_F4_53 ); 
OneRegister MUX1_F4_RO54(clk, write2_55, CompOut_F4, REGofMAX1DataOut_F4_54 ); 
OneRegister MUX1_F4_RO55(clk, write2_56, CompOut_F4, REGofMAX1DataOut_F4_55 ); 
OneRegister MUX1_F4_RO56(clk, write2_57, CompOut_F4, REGofMAX1DataOut_F4_56 ); 
OneRegister MUX1_F4_RO57(clk, write2_58, CompOut_F4, REGofMAX1DataOut_F4_57 ); 
OneRegister MUX1_F4_RO58(clk, write2_59, CompOut_F4, REGofMAX1DataOut_F4_58 ); 
OneRegister MUX1_F4_RO59(clk, write2_60, CompOut_F4, REGofMAX1DataOut_F4_59 ); 
OneRegister MUX1_F4_RO60(clk, write2_61, CompOut_F4, REGofMAX1DataOut_F4_60 ); 
OneRegister MUX1_F4_RO61(clk, write2_62, CompOut_F4, REGofMAX1DataOut_F4_61 ); 
OneRegister MUX1_F4_RO62(clk, write2_63, CompOut_F4, REGofMAX1DataOut_F4_62 ); 
OneRegister MUX1_F4_RO63(clk, write2_64, CompOut_F4, REGofMAX1DataOut_F4_63 ); 
OneRegister MUX1_F4_RO64(clk, write2_65, CompOut_F4, REGofMAX1DataOut_F4_64 ); 
OneRegister MUX1_F4_RO65(clk, write2_66, CompOut_F4, REGofMAX1DataOut_F4_65 ); 
OneRegister MUX1_F4_RO66(clk, write2_67, CompOut_F4, REGofMAX1DataOut_F4_66 ); 
OneRegister MUX1_F4_RO67(clk, write2_68, CompOut_F4, REGofMAX1DataOut_F4_67 ); 
OneRegister MUX1_F4_RO68(clk, write2_69, CompOut_F4, REGofMAX1DataOut_F4_68 ); 
OneRegister MUX1_F4_RO69(clk, write2_70, CompOut_F4, REGofMAX1DataOut_F4_69 ); 
OneRegister MUX1_F4_RO70(clk, write2_71, CompOut_F4, REGofMAX1DataOut_F4_70 ); 
OneRegister MUX1_F4_RO71(clk, write2_72, CompOut_F4, REGofMAX1DataOut_F4_71 ); 
OneRegister MUX1_F4_RO72(clk, write2_73, CompOut_F4, REGofMAX1DataOut_F4_72 ); 
OneRegister MUX1_F4_RO73(clk, write2_74, CompOut_F4, REGofMAX1DataOut_F4_73 ); 
OneRegister MUX1_F4_RO74(clk, write2_75, CompOut_F4, REGofMAX1DataOut_F4_74 ); 
OneRegister MUX1_F4_RO75(clk, write2_76, CompOut_F4, REGofMAX1DataOut_F4_75 ); 
OneRegister MUX1_F4_RO76(clk, write2_77, CompOut_F4, REGofMAX1DataOut_F4_76 ); 
OneRegister MUX1_F4_RO77(clk, write2_78, CompOut_F4, REGofMAX1DataOut_F4_77 ); 
OneRegister MUX1_F4_RO78(clk, write2_79, CompOut_F4, REGofMAX1DataOut_F4_78 ); 
OneRegister MUX1_F4_RO79(clk, write2_80, CompOut_F4, REGofMAX1DataOut_F4_79 ); 
OneRegister MUX1_F4_RO80(clk, write2_81, CompOut_F4, REGofMAX1DataOut_F4_80 ); 
OneRegister MUX1_F4_RO81(clk, write2_82, CompOut_F4, REGofMAX1DataOut_F4_81 ); 
OneRegister MUX1_F4_RO82(clk, write2_83, CompOut_F4, REGofMAX1DataOut_F4_82 ); 
OneRegister MUX1_F4_RO83(clk, write2_84, CompOut_F4, REGofMAX1DataOut_F4_83 ); 
OneRegister MUX1_F4_RO84(clk, write2_85, CompOut_F4, REGofMAX1DataOut_F4_84 ); 
OneRegister MUX1_F4_RO85(clk, write2_86, CompOut_F4, REGofMAX1DataOut_F4_85 ); 
OneRegister MUX1_F4_RO86(clk, write2_87, CompOut_F4, REGofMAX1DataOut_F4_86 ); 
OneRegister MUX1_F4_RO87(clk, write2_88, CompOut_F4, REGofMAX1DataOut_F4_87 ); 
OneRegister MUX1_F4_RO88(clk, write2_89, CompOut_F4, REGofMAX1DataOut_F4_88 ); 
OneRegister MUX1_F4_RO89(clk, write2_90, CompOut_F4, REGofMAX1DataOut_F4_89 ); 
OneRegister MUX1_F4_RO90(clk, write2_91, CompOut_F4, REGofMAX1DataOut_F4_90 ); 
OneRegister MUX1_F4_RO91(clk, write2_92, CompOut_F4, REGofMAX1DataOut_F4_91 ); 
OneRegister MUX1_F4_RO92(clk, write2_93, CompOut_F4, REGofMAX1DataOut_F4_92 ); 
OneRegister MUX1_F4_RO93(clk, write2_94, CompOut_F4, REGofMAX1DataOut_F4_93 ); 
OneRegister MUX1_F4_RO94(clk, write2_95, CompOut_F4, REGofMAX1DataOut_F4_94 ); 
OneRegister MUX1_F4_RO95(clk, write2_96, CompOut_F4, REGofMAX1DataOut_F4_95 ); 
OneRegister MUX1_F4_RO96(clk, write2_97, CompOut_F4, REGofMAX1DataOut_F4_96 ); 
OneRegister MUX1_F4_RO97(clk, write2_98, CompOut_F4, REGofMAX1DataOut_F4_97 ); 
OneRegister MUX1_F4_RO98(clk, write2_99, CompOut_F4, REGofMAX1DataOut_F4_98 ); 
OneRegister MUX1_F4_RO99(clk, write2_100, CompOut_F4, REGofMAX1DataOut_F4_99 ); 
OneRegister MUX1_F4_RO100(clk, write2_101, CompOut_F4, REGofMAX1DataOut_F4_100 ); 
OneRegister MUX1_F4_RO101(clk, write2_102, CompOut_F4, REGofMAX1DataOut_F4_101 ); 
OneRegister MUX1_F4_RO102(clk, write2_103, CompOut_F4, REGofMAX1DataOut_F4_102 ); 
OneRegister MUX1_F4_RO103(clk, write2_104, CompOut_F4, REGofMAX1DataOut_F4_103 ); 
OneRegister MUX1_F4_RO104(clk, write2_105, CompOut_F4, REGofMAX1DataOut_F4_104 ); 
OneRegister MUX1_F4_RO105(clk, write2_106, CompOut_F4, REGofMAX1DataOut_F4_105 ); 
OneRegister MUX1_F4_RO106(clk, write2_107, CompOut_F4, REGofMAX1DataOut_F4_106 ); 
OneRegister MUX1_F4_RO107(clk, write2_108, CompOut_F4, REGofMAX1DataOut_F4_107 ); 
OneRegister MUX1_F4_RO108(clk, write2_109, CompOut_F4, REGofMAX1DataOut_F4_108 ); 
OneRegister MUX1_F4_RO109(clk, write2_110, CompOut_F4, REGofMAX1DataOut_F4_109 ); 
OneRegister MUX1_F4_RO110(clk, write2_111, CompOut_F4, REGofMAX1DataOut_F4_110 ); 
OneRegister MUX1_F4_RO111(clk, write2_112, CompOut_F4, REGofMAX1DataOut_F4_111 ); 
OneRegister MUX1_F4_RO112(clk, write2_113, CompOut_F4, REGofMAX1DataOut_F4_112 ); 
OneRegister MUX1_F4_RO113(clk, write2_114, CompOut_F4, REGofMAX1DataOut_F4_113 ); 
OneRegister MUX1_F4_RO114(clk, write2_115, CompOut_F4, REGofMAX1DataOut_F4_114 ); 
OneRegister MUX1_F4_RO115(clk, write2_116, CompOut_F4, REGofMAX1DataOut_F4_115 ); 
OneRegister MUX1_F4_RO116(clk, write2_117, CompOut_F4, REGofMAX1DataOut_F4_116 ); 
OneRegister MUX1_F4_RO117(clk, write2_118, CompOut_F4, REGofMAX1DataOut_F4_117 ); 
OneRegister MUX1_F4_RO118(clk, write2_119, CompOut_F4, REGofMAX1DataOut_F4_118 ); 
OneRegister MUX1_F4_RO119(clk, write2_120, CompOut_F4, REGofMAX1DataOut_F4_119 ); 
OneRegister MUX1_F4_RO120(clk, write2_121, CompOut_F4, REGofMAX1DataOut_F4_120 ); 
OneRegister MUX1_F4_RO121(clk, write2_122, CompOut_F4, REGofMAX1DataOut_F4_121 ); 
OneRegister MUX1_F4_RO122(clk, write2_123, CompOut_F4, REGofMAX1DataOut_F4_122 ); 
OneRegister MUX1_F4_RO123(clk, write2_124, CompOut_F4, REGofMAX1DataOut_F4_123 ); 
OneRegister MUX1_F4_RO124(clk, write2_125, CompOut_F4, REGofMAX1DataOut_F4_124 ); 
OneRegister MUX1_F4_RO125(clk, write2_126, CompOut_F4, REGofMAX1DataOut_F4_125 ); 
OneRegister MUX1_F4_RO126(clk, write2_127, CompOut_F4, REGofMAX1DataOut_F4_126 ); 
OneRegister MUX1_F4_RO127(clk, write2_128, CompOut_F4, REGofMAX1DataOut_F4_127 ); 
OneRegister MUX1_F4_RO128(clk, write2_129, CompOut_F4, REGofMAX1DataOut_F4_128 ); 
OneRegister MUX1_F4_RO129(clk, write2_130, CompOut_F4, REGofMAX1DataOut_F4_129 ); 
OneRegister MUX1_F4_RO130(clk, write2_131, CompOut_F4, REGofMAX1DataOut_F4_130 ); 
OneRegister MUX1_F4_RO131(clk, write2_132, CompOut_F4, REGofMAX1DataOut_F4_131 ); 
OneRegister MUX1_F4_RO132(clk, write2_133, CompOut_F4, REGofMAX1DataOut_F4_132 ); 
OneRegister MUX1_F4_RO133(clk, write2_134, CompOut_F4, REGofMAX1DataOut_F4_133 ); 
OneRegister MUX1_F4_RO134(clk, write2_135, CompOut_F4, REGofMAX1DataOut_F4_134 ); 
OneRegister MUX1_F4_RO135(clk, write2_136, CompOut_F4, REGofMAX1DataOut_F4_135 ); 
OneRegister MUX1_F4_RO136(clk, write2_137, CompOut_F4, REGofMAX1DataOut_F4_136 ); 
OneRegister MUX1_F4_RO137(clk, write2_138, CompOut_F4, REGofMAX1DataOut_F4_137 ); 
OneRegister MUX1_F4_RO138(clk, write2_139, CompOut_F4, REGofMAX1DataOut_F4_138 ); 
OneRegister MUX1_F4_RO139(clk, write2_140, CompOut_F4, REGofMAX1DataOut_F4_139 ); 
OneRegister MUX1_F4_RO140(clk, write2_141, CompOut_F4, REGofMAX1DataOut_F4_140 ); 
OneRegister MUX1_F4_RO141(clk, write2_142, CompOut_F4, REGofMAX1DataOut_F4_141 ); 
OneRegister MUX1_F4_RO142(clk, write2_143, CompOut_F4, REGofMAX1DataOut_F4_142 ); 
OneRegister MUX1_F4_RO143(clk, write2_144, CompOut_F4, REGofMAX1DataOut_F4_143 ); 



endmodule

