module compTB();
reg clk;
reg [33:0] A , B  ;
localparam period = 100; 
wire unorderedAB,  AltB , AeqB , AgtB , AleB , AgeB ;
FPComparator_8_23_F400_uid2 CompInstanceAB (clk , A , B ,  unorderedAB,  AltB , AeqB , AgtB , AleB , AgeB );
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	
A   <=34'b0100111111110000000000000000000000;
B   <=34'b0110111111111000000000000000000000;
#period;
end 
endmodule



module maxpoolTB();
reg clk;
reg [33:0] A , B , C, D ;
localparam period = 100; 
wire [33:0] Data;
COMPARATOR_MAX_TRY_tssssst   TBinstance ( clk, A,B, C, D, Data) ;
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	
A   <=34'b0100111111110000000000000000000000; //1.5
B   <=34'b0110111111111000000000000000000000; //-1.75
C   <=34'b0100111111101000000000000000000000; //1.25
D   <=34'b0000000000000000000000000000000000; //0
#period;

end 
endmodule




module AdderTB();
reg clk;
reg [33:0] A , B ;
localparam period = 100; 
wire [33:0] C;
FPAdd_8_23_F400_uid2 AdderInstance (clk,  A ,  B ,  C  );
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	
A   <=34'b0100111111110000000000000000000000; //1.5
B   <=34'b0110111111111000000000000000000000; //-1.75

#period;
//0110111110100000000000000000000000 the answer is after 7.5 cycles
end 
endmodule


module AdderTB66bits();
reg clk;
reg [65:0] A , B ;
localparam period = 100; 
wire [65:0] C;
DoubleAdder AdderInstance (clk,  A ,  B ,  C  );
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	
A   <=66'b011011111111110100000000000000000000000000000000000000000000000000; //-1.25
B   <=66'b010011111111110100000000000000000000000000000000000000000000000000; //1.25

#period;
//000000000000000000000000000000000000000000000000000000000000000000 the answer is after 9.5 cycles
end 
endmodule


module Adder5numbersTB(); //reset = 1 flawl bs, mac start = 1, mac end = 0, change a every 13 cycles
reg clk, MAC_start, MAC_end, resetTheCounter;
reg [33:0] A ;

localparam period = 100; 
wire [33:0] Z;
AdderAcc_5 INSTANCENAME (A, clk, Z, MAC_start, MAC_end, resetTheCounter);
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	
 resetTheCounter = 1;
 MAC_start = 0;
 MAC_end = 0;
 #20;
 resetTheCounter = 0;
 MAC_start = 1;
 MAC_end = 0;

A   <=34'b0100111111110000000000000000000000; //1.5
 #1300;
A   <=34'b0110111111111000000000000000000000; //-1.75
 #1300;
A  <=34'b0100111111101000000000000000000000; //1.25
 #1300;
A  <=34'b0000000000000000000000000000000000; //0
 #1300;
A   <= 34'b0101000000011000000000000000000000; //3.5
 #1300;
 MAC_start = 0;
 MAC_end = 1;
 //0110111110100000000000000000000000   //-.25
 //0100111111100000000000000000000000   //1
 //0100111111100000000000000000000000   //1
//0101000000100100000000000000000000 //4.5
end 
endmodule



//FPMult_8_23_8_23_8_23_uid2_F400_uid3 MultiplierInstance (clk, A , B , R )

module MulTB();
reg clk;
reg [33:0] A , B  ;
localparam period = 100; 
wire [33:0] R ;
FPMult_8_23_8_23_8_23_uid2_F400_uid3 MultiplierInstance (clk, A , B , R );
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	
A   <=34'b0110111111110000000000000000000000; //-1.5
B   <=34'b0101000000000000000000000000000000; //2
#period;
//-3 //0111000000010000000000000000000000 AFTER HALF CYCLE
end 
endmodule


//

module MAC9numbersTB(); //reset = 1 flawl bs, mac start = 1, mac end = 0, change a every 13 cycles
reg clk, MAC_start, MAC_end, resetTheCounter;
reg [33:0] A, B ;

localparam period = 100; 
wire [33:0] Z;

MAC_9 macinstance (A, B, clk, Z, MAC_start, MAC_end, resetTheCounter);

always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	
 resetTheCounter = 1;
 MAC_start = 0;
 MAC_end = 0;
 #20;
 resetTheCounter = 0;
 MAC_start = 1;
 MAC_end = 0;

A   <=34'b0100111111110000000000000000000000; //1.5
B   <= 34'b0000000000000000000000000000000000; //0
 #1300;
A   <=34'b0110111111111000000000000000000000; //-1.75
B   <=34'b0110111111111000000000000000000000; //-1.75
 #1300;
A  <=34'b0100111111101000000000000000000000; //1.25
B  <=34'b0100111111101000000000000000000000; //1.25
 #1300;
A  <=34'b0000000000000000000000000000000000; //0
B   <= 34'b0101000000011000000000000000000000; //3.5
 #1300;
A   <= 34'b0101000000011000000000000000000000; //3.5
B   <=34'b0100111111110000000000000000000000; //1.5
 #1300;
A   <=34'b0110111111111000000000000000000000; //-1.75
B   <=34'b0110111111111000000000000000000000; //-1.75
 #1300;
A  <=34'b0100111111101000000000000000000000; //1.25
B  <=34'b0100111111101000000000000000000000; //1.25
 #1300;
A  <=34'b0000000000000000000000000000000000; //0
B   <= 34'b0101000000011000000000000000000000; //3.5
 #1300;
A   <= 34'b0101000000011000000000000000000000; //3.5
B   <=34'b0110111111110000000000000000000000; //-1.5
 #1300;
 MAC_start = 0;
 MAC_end = 1;
 //0101000001000101000000000000000000   //9.25

end 
endmodule



module L2toL4TB();
reg clk, Conv2LayerStart;
wire MAX2LayerFinish;


reg [33:0] REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143  ;

wire [33:0] MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 ;


localparam period = 100; 



MERGEHOPE_L3_L4  L2toL4instance (clk, Conv2LayerStart, MAX2LayerFinish
,REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143 
,MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 
 );
 
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	
Conv2LayerStart <= 1'b1;


REGofMAX1DataOut_F1_0 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_1 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_2 <= 34'b0101000010001001001010011000100100   ;
REGofMAX1DataOut_F1_3 <= 34'b0101000011011010101110111010101011   ;
REGofMAX1DataOut_F1_4 <= 34'b0101000011101101011100011010011001   ;
REGofMAX1DataOut_F1_5 <= 34'b0101000011110111111001101110011100   ;
REGofMAX1DataOut_F1_6 <= 34'b0101000011111011111110111101111101   ;
REGofMAX1DataOut_F1_7 <= 34'b0101000011100100110011001010100100   ;
REGofMAX1DataOut_F1_8 <= 34'b0101000010100001110100011111010101   ;
REGofMAX1DataOut_F1_9 <= 34'b0101000000011000100011010010011010   ;
REGofMAX1DataOut_F1_10 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_11 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_12 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_13 <= 34'b0101000010000010010100101011111100   ;
REGofMAX1DataOut_F1_14 <= 34'b0101000011100100011000110011101011   ;
REGofMAX1DataOut_F1_15 <= 34'b0101000100000000001110000111010010   ;
REGofMAX1DataOut_F1_16 <= 34'b0101000100000101100100100101111011   ;
REGofMAX1DataOut_F1_17 <= 34'b0101000100001010001111000011111110   ;
REGofMAX1DataOut_F1_18 <= 34'b0101000100001100010110010100101011   ;
REGofMAX1DataOut_F1_19 <= 34'b0101000100001100001110101111000110   ;
REGofMAX1DataOut_F1_20 <= 34'b0101000100000100110010111001011111   ;
REGofMAX1DataOut_F1_21 <= 34'b0101000011001011110101100000000001   ;
REGofMAX1DataOut_F1_22 <= 34'b0101000001011111001100001000100011   ;
REGofMAX1DataOut_F1_23 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_24 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_25 <= 34'b0101000011010011001111111100000010   ;
REGofMAX1DataOut_F1_26 <= 34'b0101000011100110100000000000011000   ;
REGofMAX1DataOut_F1_27 <= 34'b0101000011110100010101011011111111   ;
REGofMAX1DataOut_F1_28 <= 34'b0101000011110101110000101000011001   ;
REGofMAX1DataOut_F1_29 <= 34'b0101000011010100001001111111101101   ;
REGofMAX1DataOut_F1_30 <= 34'b0101000011101111100100110011110010   ;
REGofMAX1DataOut_F1_31 <= 34'b0101000100000111100100011110100010   ;
REGofMAX1DataOut_F1_32 <= 34'b0101000100001001110101001001000010   ;
REGofMAX1DataOut_F1_33 <= 34'b0101000011111111100011110100101001   ;
REGofMAX1DataOut_F1_34 <= 34'b0101000011001010110010011101010100   ;
REGofMAX1DataOut_F1_35 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_36 <= 34'b0101000001101000001000000001011001   ;
REGofMAX1DataOut_F1_37 <= 34'b0101000011010000100000111101000000   ;
REGofMAX1DataOut_F1_38 <= 34'b0101000011011011001111100111100010   ;
REGofMAX1DataOut_F1_39 <= 34'b0101000010110110100111110100000111   ;
REGofMAX1DataOut_F1_40 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_41 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_42 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_43 <= 34'b0101000001010111111111011101011101   ;
REGofMAX1DataOut_F1_44 <= 34'b0101000011111101011000011111011100   ;
REGofMAX1DataOut_F1_45 <= 34'b0101000011111111101110010010101000   ;
REGofMAX1DataOut_F1_46 <= 34'b0101000011101001110000101001100111   ;
REGofMAX1DataOut_F1_47 <= 34'b0101000010000101101110111111110100   ;
REGofMAX1DataOut_F1_48 <= 34'b0101000010001101000111011001001110   ;
REGofMAX1DataOut_F1_49 <= 34'b0101000011000001001101000100101111   ;
REGofMAX1DataOut_F1_50 <= 34'b0101000011001000001000110010100111   ;
REGofMAX1DataOut_F1_51 <= 34'b0101000010101110110110101011110110   ;
REGofMAX1DataOut_F1_52 <= 34'b0101000001010000111101001010010100   ;
REGofMAX1DataOut_F1_53 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_54 <= 34'b0101000000111100111111110101000000   ;
REGofMAX1DataOut_F1_55 <= 34'b0000000000000000000000000000000000   ;
REGofMAX1DataOut_F1_56 <= 34'b0101000010110010100011110000111000   ;
REGofMAX1DataOut_F1_57 <= 34'b0101000011101111011110111111000011   ;
REGofMAX1DataOut_F1_58 <= 34'b0101000011101101100011000001111000   ;
REGofMAX1DataOut_F1_59 <= 34'b0101000010110111011110011011101110   ;
REGofMAX1DataOut_F1_60 <= 34'b0101000010111111010010110011100101   ;
REGofMAX1DataOut_F1_61 <= 34'b0101000011000111100111011100101110   ;
REGofMAX1DataOut_F1_62 <= 34'b0101000011001100110100010100001111   ;
REGofMAX1DataOut_F1_63 <= 34'b0101000011011000110010001100011100   ;
REGofMAX1DataOut_F1_64 <= 34'b0101000011001100110111001111111110 ;
REGofMAX1DataOut_F1_65 <= 34'b0101000000111111110001010001010101 ;
REGofMAX1DataOut_F1_66 <= 34'b0000000000000000000000000000000000 ;
REGofMAX1DataOut_F1_67 <= 34'b0000000000000000000000000000000000 ;
REGofMAX1DataOut_F1_68 <= 34'b0000000000000000000000000000000000 ;
REGofMAX1DataOut_F1_69 <= 34'b0101000011100010100111100110111100 ;
REGofMAX1DataOut_F1_70 <= 34'b0101000011100111001000001101000010 ;
REGofMAX1DataOut_F1_71 <= 34'b0101000011001110101001011111100000  ;
REGofMAX1DataOut_F1_72 <= 34'b0101000010100010101011000011111111  ;
REGofMAX1DataOut_F1_73 <= 34'b0101000011000101101010000100010101  ;
REGofMAX1DataOut_F1_74 <= 34'b0101000011100011001011111100001110  ;
REGofMAX1DataOut_F1_75 <= 34'b0101000011101000010111011010011111  ;
REGofMAX1DataOut_F1_76 <= 34'b0101000011010100010010000110011111  ;
REGofMAX1DataOut_F1_77 <= 34'b0100111111100111110001110000100011  ;
REGofMAX1DataOut_F1_78 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F1_79 <= 34'b0101000010011001011000110111000110  ;
REGofMAX1DataOut_F1_80 <= 34'b0101000010010110011111000110101100  ;
REGofMAX1DataOut_F1_81 <= 34'b0101000011000111000011100011100011  ;
REGofMAX1DataOut_F1_82 <= 34'b0101000011100010010111011101010110  ;
REGofMAX1DataOut_F1_83 <= 34'b0101000011001111100011100111001111  ;
REGofMAX1DataOut_F1_84 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F1_85 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F1_86 <= 34'b0101000011100100101011110011010010  ;
REGofMAX1DataOut_F1_87 <= 34'b0101000100000100000011111000001110  ;
REGofMAX1DataOut_F1_88 <= 34'b0101000100000010001100110000001110  ;
REGofMAX1DataOut_F1_89 <= 34'b0101000011001011010011101101001011  ;
REGofMAX1DataOut_F1_90 <= 34'b0101000011000000110111001101100101  ;
REGofMAX1DataOut_F1_91 <= 34'b0101000011100101011111101000110011  ;
REGofMAX1DataOut_F1_92 <= 34'b0101000011100010101110100011011001  ;
REGofMAX1DataOut_F1_93 <= 34'b0101000010100011110001111000100010  ;
REGofMAX1DataOut_F1_94 <= 34'b0101000011000110101110100111000011  ;
REGofMAX1DataOut_F1_95 <= 34'b0101000011000010001011110000110010  ;
REGofMAX1DataOut_F1_96 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F1_97 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F1_98 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F1_99 <= 34'b0101000100000010111100001100001101  ;
REGofMAX1DataOut_F1_100 <= 34'b0101000100001011000010110010010011   ;
REGofMAX1DataOut_F1_101 <= 34'b0101000100001100011101110101110110  ;
REGofMAX1DataOut_F1_102 <= 34'b0101000100001001010001101100111000  ;
REGofMAX1DataOut_F1_103 <= 34'b0101000100000011100011010100101011  ;
REGofMAX1DataOut_F1_104 <= 34'b0101000011110001110101100110010000  ;
REGofMAX1DataOut_F1_105 <= 34'b0101000010110000000100000101101011  ;
REGofMAX1DataOut_F1_106 <= 34'b0101000010100011110101101111101010  ;
REGofMAX1DataOut_F1_107 <= 34'b0101000010000000011110010100000110  ;
REGofMAX1DataOut_F1_108 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F1_109 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_110 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_111 <= 34'b0101000010100101101101011111101010  ; 
REGofMAX1DataOut_F1_112 <= 34'b0101000100000010000010000010000110  ; 
REGofMAX1DataOut_F1_113 <= 34'b0101000100001011100001001010110100  ; 
REGofMAX1DataOut_F1_114 <= 34'b0101000100001011001100100110010000  ; 
REGofMAX1DataOut_F1_115 <= 34'b0101000100000001111100101100101000  ; 
REGofMAX1DataOut_F1_116 <= 34'b0101000010110001011010001000101000  ; 
REGofMAX1DataOut_F1_117 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_118 <= 34'b0101000010010000100111010000010100  ; 
REGofMAX1DataOut_F1_119 <= 34'b0101000000011001111000001011011111  ; 
REGofMAX1DataOut_F1_120 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F1_121 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_122 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_123 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_124 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_125 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_126 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_127 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_128 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_129 <= 34'b0101000001001101101100011111100011  ; 
REGofMAX1DataOut_F1_130 <= 34'b0101000001010100100001101010100011  ; 
REGofMAX1DataOut_F1_131 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_132 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_133 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_134 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_135 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_136 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_137 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_138 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_139 <= 34'b0101000000000100100101001000000110  ; 
REGofMAX1DataOut_F1_140 <= 34'b0101000001001000111111101110011010  ; 
REGofMAX1DataOut_F1_141 <= 34'b0101000001100110101000010110101111  ; 
REGofMAX1DataOut_F1_142 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F1_143 <= 34'b0000000000000000000000000000000000  ; 


REGofMAX1DataOut_F2_0 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_1 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_2 <= 34'b0101000001101001000011101000011100  ;
REGofMAX1DataOut_F2_3 <= 34'b0101000011001101110000111010110100  ;
REGofMAX1DataOut_F2_4 <= 34'b0101000011101000011101110000001000  ;
REGofMAX1DataOut_F2_5 <= 34'b0101000011101101001110100111001000  ;
REGofMAX1DataOut_F2_6 <= 34'b0101000011101011111010011111111000  ;
REGofMAX1DataOut_F2_7 <= 34'b0101000011100000101101110001001111  ;
REGofMAX1DataOut_F2_8 <= 34'b0101000010011111100010000011111010  ;
REGofMAX1DataOut_F2_9 <= 34'b0100111100110100100000011101011111  ;
REGofMAX1DataOut_F2_10 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_11 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_12 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_13 <= 34'b0101000001001011111010111110100010  ;
REGofMAX1DataOut_F2_14 <= 34'b0101000010111010101101000101101111  ;
REGofMAX1DataOut_F2_15 <= 34'b0101000011100010011000001101000001  ;
REGofMAX1DataOut_F2_16 <= 34'b0101000011011101100001000111110010  ;
REGofMAX1DataOut_F2_17 <= 34'b0101000011000101111010000101100110  ;
REGofMAX1DataOut_F2_18 <= 34'b0101000011100101011000000011100000  ;
REGofMAX1DataOut_F2_19 <= 34'b0101000011101110000001001111010100  ;
REGofMAX1DataOut_F2_20 <= 34'b0101000011101101111011000100111111  ;
REGofMAX1DataOut_F2_21 <= 34'b0101000011000101100100110010100100  ;
REGofMAX1DataOut_F2_22 <= 34'b0100111111101011101111100010011100  ;
REGofMAX1DataOut_F2_23 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_24 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_25 <= 34'b0101000010011111110011110000000101  ;
REGofMAX1DataOut_F2_26 <= 34'b0101000001101111010011100001100111  ;
REGofMAX1DataOut_F2_27 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_28 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_29 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_30 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_31 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_32 <= 34'b0101000011101001011111000111001000  ;
REGofMAX1DataOut_F2_33 <= 34'b0101000011100100101101001010101000  ;
REGofMAX1DataOut_F2_34 <= 34'b0101000010110100011110111111011000  ;
REGofMAX1DataOut_F2_35 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_36 <= 34'b0101000001000000100101011110100111  ;
REGofMAX1DataOut_F2_37 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_38 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_39 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_40 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_41 <= 34'b0101000010111101011000100100001110  ;
REGofMAX1DataOut_F2_42 <= 34'b0101000011000001101100010010011100  ;
REGofMAX1DataOut_F2_43 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_44 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_45 <= 34'b0101000011010001010110010111011111  ;
REGofMAX1DataOut_F2_46 <= 34'b0101000011001111010101100100011100  ;
REGofMAX1DataOut_F2_47 <= 34'b0101000000110011001100000101001111  ;
REGofMAX1DataOut_F2_48 <= 34'b0101000001000010011110111001011010  ;
REGofMAX1DataOut_F2_49 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_50 <= 34'b0101000010100110011101000111100111  ;
REGofMAX1DataOut_F2_51 <= 34'b0101000011010100000010101111101110  ;
REGofMAX1DataOut_F2_52 <= 34'b0101000011001111100000111000111101  ;
REGofMAX1DataOut_F2_53 <= 34'b0101000010101101011001000110010100  ;
REGofMAX1DataOut_F2_54 <= 34'b0101000011010100001001011101011111  ;
REGofMAX1DataOut_F2_55 <= 34'b0101000010111011101010111000101000  ;
REGofMAX1DataOut_F2_56 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_57 <= 34'b0101000010000010100101110110000001  ;
REGofMAX1DataOut_F2_58 <= 34'b0101000010111001110000001001000010  ;
REGofMAX1DataOut_F2_59 <= 34'b0101000010001001111011111110101111  ;
REGofMAX1DataOut_F2_60 <= 34'b0101000001011110101011000000100010  ;
REGofMAX1DataOut_F2_61 <= 34'b0101000010101101000011100111101011  ;
REGofMAX1DataOut_F2_62 <= 34'b0101000010101100001101000110111110  ;
REGofMAX1DataOut_F2_63 <= 34'b0101000010101011111101011110101000  ;
REGofMAX1DataOut_F2_64 <= 34'b0101000010001011010100111000010001  ;
REGofMAX1DataOut_F2_65 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_66 <= 34'b0101000010100010100101101000101000  ;
REGofMAX1DataOut_F2_67 <= 34'b0101000011001100011001011011101000  ;
REGofMAX1DataOut_F2_68 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_69 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_70 <= 34'b0101000010110110011101110010110000  ;
REGofMAX1DataOut_F2_71 <= 34'b0101000010010000010000101000000000  ;
REGofMAX1DataOut_F2_72 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_73 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_74 <= 34'b0101000001101010110011001011001011  ;
REGofMAX1DataOut_F2_75 <= 34'b0101000010110101101001101111000001  ;
REGofMAX1DataOut_F2_76 <= 34'b0101000010110100111111000010100110  ;
REGofMAX1DataOut_F2_77 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_78 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_79 <= 34'b0101000010110000111000111101001011  ;
REGofMAX1DataOut_F2_80 <= 34'b0101000010111011100001110100001100  ;
REGofMAX1DataOut_F2_81 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_82 <= 34'b0101000010010101010010010000000010  ;
REGofMAX1DataOut_F2_83 <= 34'b0101000010010100011101101000110101  ;
REGofMAX1DataOut_F2_84 <= 34'b0101000010101001010101000110110110  ;
REGofMAX1DataOut_F2_85 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_86 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_87 <= 34'b0101000011010111101000010101101000  ;
REGofMAX1DataOut_F2_88 <= 34'b0101000011100110010100001100110110  ;
REGofMAX1DataOut_F2_89 <= 34'b0101000011000001111011000011010011  ;
REGofMAX1DataOut_F2_90 <= 34'b0101000010100111111110110100101110  ;
REGofMAX1DataOut_F2_91 <= 34'b0101000011000010101010011101101111  ;
REGofMAX1DataOut_F2_92 <= 34'b0101000011001101111011010101010000  ;
REGofMAX1DataOut_F2_93 <= 34'b0101000010001010111110010101111011  ;
REGofMAX1DataOut_F2_94 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_95 <= 34'b0101000001100110010001111000001000  ;
REGofMAX1DataOut_F2_96 <= 34'b0101000010100101010010000000100000  ;
REGofMAX1DataOut_F2_97 <= 34'b0101000011000000001111100001100100  ;
REGofMAX1DataOut_F2_98 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_99 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_100 <= 34'b0101000011101110000010010111101000  ;
REGofMAX1DataOut_F2_101 <= 34'b0101000011110001011010100001000011  ;
REGofMAX1DataOut_F2_102 <= 34'b0101000011101001010111011111011001  ;
REGofMAX1DataOut_F2_103 <= 34'b0101000011011000111110110111010010  ;
REGofMAX1DataOut_F2_104 <= 34'b0101000010010000101001100110011110  ;
REGofMAX1DataOut_F2_105 <= 34'b0101000010011110010111111110010001  ;
REGofMAX1DataOut_F2_106 <= 34'b0100111111101010001111000010011100  ;
REGofMAX1DataOut_F2_107 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_108 <= 34'b0101000001000000010100100001101101  ;
REGofMAX1DataOut_F2_109 <= 34'b0101000011000110001010101011000101  ; 
REGofMAX1DataOut_F2_110 <= 34'b0101000011000011001101011010110110  ; 
REGofMAX1DataOut_F2_111 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_112 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_113 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_114 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_115 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_116 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_117 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_118 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_119 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_120 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F2_121 <= 34'b0101000010001110011101111100011010  ; 
REGofMAX1DataOut_F2_122 <= 34'b0101000011001010000010101101001111  ; 
REGofMAX1DataOut_F2_123 <= 34'b0101000011000100110010010000001110  ; 
REGofMAX1DataOut_F2_124 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_125 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_126 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_127 <= 34'b0101000001110001010010111001100001  ; 
REGofMAX1DataOut_F2_128 <= 34'b0101000010001111100100011100110110  ; 
REGofMAX1DataOut_F2_129 <= 34'b0101000001101011111001001010111010  ; 
REGofMAX1DataOut_F2_130 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_131 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_132 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_133 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_134 <= 34'b0101000010110011111101110100101000  ; 
REGofMAX1DataOut_F2_135 <= 34'b0101000011100001110000001111111000  ; 
REGofMAX1DataOut_F2_136 <= 34'b0101000011100101010101001010011000  ; 
REGofMAX1DataOut_F2_137 <= 34'b0101000011100111101101100010000001  ; 
REGofMAX1DataOut_F2_138 <= 34'b0101000011010111001011100001010010  ; 
REGofMAX1DataOut_F2_139 <= 34'b0101000011001111101011000100000010  ; 
REGofMAX1DataOut_F2_140 <= 34'b0101000010011010001110100110001101  ; 
REGofMAX1DataOut_F2_141 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_142 <= 34'b0000000000000000000000000000000000  ; 
REGofMAX1DataOut_F2_143 <= 34'b0000000000000000000000000000000000  ; 


REGofMAX1DataOut_F3_0 <= 34'b0100111011001110110001011100111001  ;
REGofMAX1DataOut_F3_1 <= 34'b0100111011001110110001011100111001  ;
REGofMAX1DataOut_F3_2 <= 34'b0101000010000010011111001100000110  ;
REGofMAX1DataOut_F3_3 <= 34'b0101000011001111011001000111010101  ;
REGofMAX1DataOut_F3_4 <= 34'b0101000011100111011000110101111001  ;
REGofMAX1DataOut_F3_5 <= 34'b0101000011101100011011000100001011  ;
REGofMAX1DataOut_F3_6 <= 34'b0101000011101001111000101111100011  ;
REGofMAX1DataOut_F3_7 <= 34'b0101000011000100010100111110000100  ;
REGofMAX1DataOut_F3_8 <= 34'b0101000000001110001001000101011001  ;
REGofMAX1DataOut_F3_9 <= 34'b0100111011001110110001011100111001  ;
REGofMAX1DataOut_F3_10 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_11 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_12 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_13 <= 34'b0101000001111100111111000110111111 ;
REGofMAX1DataOut_F3_14 <= 34'b0101000011101100010101100100011011 ;
REGofMAX1DataOut_F3_15 <= 34'b0101000100000011111111010100010110 ;
REGofMAX1DataOut_F3_16 <= 34'b0101000100010001110111111011011111 ;
REGofMAX1DataOut_F3_17 <= 34'b0101000100011110011111000000001011 ;
REGofMAX1DataOut_F3_18 <= 34'b0101000100100010111011010010001001 ;
REGofMAX1DataOut_F3_19 <= 34'b0101000100100000111000100111101011 ;
REGofMAX1DataOut_F3_20 <= 34'b0101000100000011111001101011001111 ;
REGofMAX1DataOut_F3_21 <= 34'b0101000010101001111111001001010101 ;
REGofMAX1DataOut_F3_22 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_23 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_24 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_25 <= 34'b0101000011011011101011101110001100 ;
REGofMAX1DataOut_F3_26 <= 34'b0101000011110101000101010110100100 ;
REGofMAX1DataOut_F3_27 <= 34'b0101000100001101010011110010011101 ;
REGofMAX1DataOut_F3_28 <= 34'b0101000100100001101010101110100011 ;
REGofMAX1DataOut_F3_29 <= 34'b0101000100100100000010000101010101 ;
REGofMAX1DataOut_F3_30 <= 34'b0101000100101010011100011010100100 ;
REGofMAX1DataOut_F3_31 <= 34'b0101000100101101110001100001000000 ;
REGofMAX1DataOut_F3_32 <= 34'b0101000100101101100111000001111110 ;
REGofMAX1DataOut_F3_33 <= 34'b0101000100001111010000010000011001 ;
REGofMAX1DataOut_F3_34 <= 34'b0101000010111011011111011011101000 ;
REGofMAX1DataOut_F3_35 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_36 <= 34'b0101000001100010000101010100100010 ;
REGofMAX1DataOut_F3_37 <= 34'b0101000011100111000101011010101001 ;
REGofMAX1DataOut_F3_38 <= 34'b0101000011110100111010000011000110 ;
REGofMAX1DataOut_F3_39 <= 34'b0101000100010010111100000011001011 ;
REGofMAX1DataOut_F3_40 <= 34'b0101000100011101100010010001010001 ;
REGofMAX1DataOut_F3_41 <= 34'b0101000100010100010100110010001011 ;
REGofMAX1DataOut_F3_42 <= 34'b0101000100001100001010111010000011 ;
REGofMAX1DataOut_F3_43 <= 34'b0101000100100101110101001110100001 ;
REGofMAX1DataOut_F3_44 <= 34'b0101000100101101001101100010111110 ;
REGofMAX1DataOut_F3_45 <= 34'b0101000100101011100010011000011001 ;
REGofMAX1DataOut_F3_46 <= 34'b0101000100000100100100100100010011 ;
REGofMAX1DataOut_F3_47 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_48 <= 34'b0101000010011000111101010110000010 ;
REGofMAX1DataOut_F3_49 <= 34'b0101000011011100110011000100110101 ;
REGofMAX1DataOut_F3_50 <= 34'b0101000100001001100101000110111110 ;
REGofMAX1DataOut_F3_51 <= 34'b0101000100011001011000111100110100 ;
REGofMAX1DataOut_F3_52 <= 34'b0101000100000111010001000100110010 ;
REGofMAX1DataOut_F3_53 <= 34'b0101000011111011010011110110001110 ;
REGofMAX1DataOut_F3_54 <= 34'b0101000011000011101101111111110000 ;
REGofMAX1DataOut_F3_55 <= 34'b0101000011101001111011001010010111 ;
REGofMAX1DataOut_F3_56 <= 34'b0101000100100100111111111001101101 ;
REGofMAX1DataOut_F3_57 <= 34'b0101000100101011100100100111011111 ;
REGofMAX1DataOut_F3_58 <= 34'b0101000100011100010001110011011011 ;
REGofMAX1DataOut_F3_59 <= 34'b0101000010111110101100000000001010 ;
REGofMAX1DataOut_F3_60 <= 34'b0101000011000100010011000001001000 ;
REGofMAX1DataOut_F3_61 <= 34'b0101000011100001110010000101011110 ;
REGofMAX1DataOut_F3_62 <= 34'b0101000100011100111010010100011101 ;
REGofMAX1DataOut_F3_63 <= 34'b0101000100100011010111011110111011 ;
REGofMAX1DataOut_F3_64 <= 34'b0101000011111000110110101000110101 ;
REGofMAX1DataOut_F3_65 <= 34'b0101000001101100111111100001010101 ;
REGofMAX1DataOut_F3_66 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_67 <= 34'b0000000000000000000000000000000000 ;
REGofMAX1DataOut_F3_68 <= 34'b0101000100000101111001110010000000 ;
REGofMAX1DataOut_F3_69 <= 34'b0101000100101000001010111001000001 ;
REGofMAX1DataOut_F3_70 <= 34'b0101000100100010111000011011011001 ;
REGofMAX1DataOut_F3_71 <= 34'b0101000011100100000110001000111010 ;
REGofMAX1DataOut_F3_72 <= 34'b0101000011000100111110000001001111 ;
REGofMAX1DataOut_F3_73 <= 34'b0101000011101100110010011100001111 ;
REGofMAX1DataOut_F3_74 <= 34'b0101000100100111000011000010110111 ;
REGofMAX1DataOut_F3_75 <= 34'b0101000100100101111001000001110101 ;
REGofMAX1DataOut_F3_76 <= 34'b0101000011110110000011100000000111 ;
REGofMAX1DataOut_F3_77 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_78 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_79 <= 34'b0101000001110100111110110101000011 ;
REGofMAX1DataOut_F3_80 <= 34'b0101000011100000001101000100111001 ;
REGofMAX1DataOut_F3_81 <= 34'b0101000100100010110100101101111110 ;
REGofMAX1DataOut_F3_82 <= 34'b0101000100100011101110111000111001 ;
REGofMAX1DataOut_F3_83 <= 34'b0101000011110100111011000000110111 ;
REGofMAX1DataOut_F3_84 <= 34'b0000000000000000000000000000000000 ;
REGofMAX1DataOut_F3_85 <= 34'b0101000011100110100100010110010110 ;
REGofMAX1DataOut_F3_86 <= 34'b0101000100101001010010010111001001 ;
REGofMAX1DataOut_F3_87 <= 34'b0101000100101110100011100010110000 ;
REGofMAX1DataOut_F3_88 <= 34'b0101000100010001100100010111000010 ;
REGofMAX1DataOut_F3_89 <= 34'b0101000010101010110110011100000011 ;
REGofMAX1DataOut_F3_90 <= 34'b0101000010101111101011001110110100 ;
REGofMAX1DataOut_F3_91 <= 34'b0101000011101011111111010110111011 ;
REGofMAX1DataOut_F3_92 <= 34'b0101000011101001000000001000100101 ;
REGofMAX1DataOut_F3_93 <= 34'b0101000100010011010011010011110110 ;
REGofMAX1DataOut_F3_94 <= 34'b0101000100100010010110100010101010 ;
REGofMAX1DataOut_F3_95 <= 34'b0101000011110100111011000010100001 ;
REGofMAX1DataOut_F3_96 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_97 <= 34'b0000000000000000000000000000000000 ;
REGofMAX1DataOut_F3_98 <= 34'b0101000100011110000101011101111101 ;
REGofMAX1DataOut_F3_99 <= 34'b0101000100101110100001010100010011 ;
REGofMAX1DataOut_F3_100 <= 34'b0101000100101101110110111000010110 ;
REGofMAX1DataOut_F3_101 <= 34'b0101000100011100000101011100111000 ;
REGofMAX1DataOut_F3_102 <= 34'b0101000100000111110000101100100110 ;
REGofMAX1DataOut_F3_103 <= 34'b0101000100000100110010110000110110 ;
REGofMAX1DataOut_F3_104 <= 34'b0101000100001000010011111011101101 ;
REGofMAX1DataOut_F3_105 <= 34'b0101000100011110100010101101101001 ;
REGofMAX1DataOut_F3_106 <= 34'b0101000100011010000010111010000000 ;
REGofMAX1DataOut_F3_107 <= 34'b0101000011010011111010010110101111 ;
REGofMAX1DataOut_F3_108 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_109 <= 34'b0000000000000000000000000000000000 ; 
REGofMAX1DataOut_F3_110 <= 34'b0101000011011100010010010100010001 ; 
REGofMAX1DataOut_F3_111 <= 34'b0101000100100101000110100111101100 ; 
REGofMAX1DataOut_F3_112 <= 34'b0101000100101110101010010001110110 ; 
REGofMAX1DataOut_F3_113 <= 34'b0101000100101011011000000101001100 ; 
REGofMAX1DataOut_F3_114 <= 34'b0101000100100100101011111011100010 ; 
REGofMAX1DataOut_F3_115 <= 34'b0101000100011001110010010110010010 ; 
REGofMAX1DataOut_F3_116 <= 34'b0101000100010111110011101101100100 ; 
REGofMAX1DataOut_F3_117 <= 34'b0101000100011011101011111010011010 ; 
REGofMAX1DataOut_F3_118 <= 34'b0101000100001010010000010001001110 ; 
REGofMAX1DataOut_F3_119 <= 34'b0101000001001001101001000001100010 ; 
REGofMAX1DataOut_F3_120 <= 34'b0100111011001110110001011100111001 ;
REGofMAX1DataOut_F3_121 <= 34'b0100111011001110110001011100111001 ; 
REGofMAX1DataOut_F3_122 <= 34'b0000000000000000000000000000000000 ; 
REGofMAX1DataOut_F3_123 <= 34'b0101000011011110010001010010011111 ; 
REGofMAX1DataOut_F3_124 <= 34'b0101000100011100001010110010110010 ; 
REGofMAX1DataOut_F3_125 <= 34'b0101000100100010100011101000110100 ; 
REGofMAX1DataOut_F3_126 <= 34'b0101000100100010000110000101100001 ; 
REGofMAX1DataOut_F3_127 <= 34'b0101000100011000001110101010001010 ; 
REGofMAX1DataOut_F3_128 <= 34'b0101000100010010000011001100110001 ; 
REGofMAX1DataOut_F3_129 <= 34'b0101000100001011111111100100111110 ; 
REGofMAX1DataOut_F3_130 <= 34'b0101000011010001000110010000111000 ; 
REGofMAX1DataOut_F3_131 <= 34'b0100111011001110110001011100111001 ; 
REGofMAX1DataOut_F3_132 <= 34'b0100111011001110110001011100111001 ; 
REGofMAX1DataOut_F3_133 <= 34'b0100111011001110110001011100111001 ; 
REGofMAX1DataOut_F3_134 <= 34'b0100111011001110110001011100111001 ; 
REGofMAX1DataOut_F3_135 <= 34'b0000000000000000000000000000000000 ; 
REGofMAX1DataOut_F3_136 <= 34'b0101000010001001101101010100011110 ; 
REGofMAX1DataOut_F3_137 <= 34'b0101000011100101101001101011101011 ; 
REGofMAX1DataOut_F3_138 <= 34'b0101000011111010111110111111101000 ; 
REGofMAX1DataOut_F3_139 <= 34'b0101000011111010101000101001000001 ; 
REGofMAX1DataOut_F3_140 <= 34'b0101000011101001010001000000011110 ; 
REGofMAX1DataOut_F3_141 <= 34'b0101000011000000100011101111001000 ; 
REGofMAX1DataOut_F3_142 <= 34'b0100111011001110110001011100111001 ; 
REGofMAX1DataOut_F3_143 <= 34'b0100111011001110110001011100111001 ; 


REGofMAX1DataOut_F4_0 <= 34'b0100111001011001000100111110011001 ;
REGofMAX1DataOut_F4_1 <= 34'b0100111001011001000100111110011001 ;
REGofMAX1DataOut_F4_2 <= 34'b0101000010011011001001100000101010 ;
REGofMAX1DataOut_F4_3 <= 34'b0101000011100110100101100100111000 ;
REGofMAX1DataOut_F4_4 <= 34'b0101000011111010000100110000111100 ;
REGofMAX1DataOut_F4_5 <= 34'b0101000011111110010001110000010110 ;
REGofMAX1DataOut_F4_6 <= 34'b0101000011101100111111011011000111 ;
REGofMAX1DataOut_F4_7 <= 34'b0101000010101000011011000011111000 ;
REGofMAX1DataOut_F4_8 <= 34'b0000000000000000000000000000000000 ;
REGofMAX1DataOut_F4_9 <= 34'b0100111001011001000100111110011001 ;
REGofMAX1DataOut_F4_10 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_11 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_12 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_13 <= 34'b0101000010010101000100110000011111  ;
REGofMAX1DataOut_F4_14 <= 34'b0101000100000000000010100011110011  ;
REGofMAX1DataOut_F4_15 <= 34'b0101000100010000011101000001010001  ;
REGofMAX1DataOut_F4_16 <= 34'b0101000100001111000100011000110111  ;
REGofMAX1DataOut_F4_17 <= 34'b0101000100001100011000000101000111  ;
REGofMAX1DataOut_F4_18 <= 34'b0101000100000111011101011110101010  ;
REGofMAX1DataOut_F4_19 <= 34'b0101000011110111100010100001110000  ;
REGofMAX1DataOut_F4_20 <= 34'b0101000010111000101111010011111100  ;
REGofMAX1DataOut_F4_21 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F4_22 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_23 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_24 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_25 <= 34'b0101000011110000000000111010010010  ;
REGofMAX1DataOut_F4_26 <= 34'b0101000100011000111010110110000010  ;
REGofMAX1DataOut_F4_27 <= 34'b0101000100011101010011011001100100  ;
REGofMAX1DataOut_F4_28 <= 34'b0101000100010101000101111111100001  ;
REGofMAX1DataOut_F4_29 <= 34'b0101000100001010000010001000110010  ;
REGofMAX1DataOut_F4_30 <= 34'b0101000100001111110100001010101010  ;
REGofMAX1DataOut_F4_31 <= 34'b0101000100010100011000110000001111  ;
REGofMAX1DataOut_F4_32 <= 34'b0101000100000110010111000001001101  ;
REGofMAX1DataOut_F4_33 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F4_34 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F4_35 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_36 <= 34'b0101000001111011011110101011110100  ;
REGofMAX1DataOut_F4_37 <= 34'b0101000100001100101111010010111111  ;
REGofMAX1DataOut_F4_38 <= 34'b0101000100011101000100101111000000  ;
REGofMAX1DataOut_F4_39 <= 34'b0101000100010010010011100100101101  ;
REGofMAX1DataOut_F4_40 <= 34'b0101000100000000011001111110011110  ;
REGofMAX1DataOut_F4_41 <= 34'b0101000011101001110000000001100111  ;
REGofMAX1DataOut_F4_42 <= 34'b0101000100001010100101000100101110  ;
REGofMAX1DataOut_F4_43 <= 34'b0101000100011101101001001010010100  ;
REGofMAX1DataOut_F4_44 <= 34'b0101000100011111101011011100110110  ;
REGofMAX1DataOut_F4_45 <= 34'b0101000011110101011010010001100000  ;
REGofMAX1DataOut_F4_46 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F4_47 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_48 <= 34'b0101000010110000100101001110010001  ;
REGofMAX1DataOut_F4_49 <= 34'b0101000100011000000001100011111100  ;
REGofMAX1DataOut_F4_50 <= 34'b0101000100100000101111111100101101  ;
REGofMAX1DataOut_F4_51 <= 34'b0101000011101101011110010010101000  ;
REGofMAX1DataOut_F4_52 <= 34'b0101000011000101011100001101110110  ;
REGofMAX1DataOut_F4_53 <= 34'b0101000011000101110000001011101100  ;
REGofMAX1DataOut_F4_54 <= 34'b0101000011100101000110010100110010  ;
REGofMAX1DataOut_F4_55 <= 34'b0101000100010111011100101011110000  ;
REGofMAX1DataOut_F4_56 <= 34'b0101000100100010000010100011001001  ;
REGofMAX1DataOut_F4_57 <= 34'b0101000100010010111101100111111011  ;
REGofMAX1DataOut_F4_58 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F4_59 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_60 <= 34'b0101000011101101100101101111101010  ;
REGofMAX1DataOut_F4_61 <= 34'b0101000100011111011111000101001101  ;
REGofMAX1DataOut_F4_62 <= 34'b0101000100100010101110010100011110  ;
REGofMAX1DataOut_F4_63 <= 34'b0101000010110111101101100000010000  ;
REGofMAX1DataOut_F4_64 <= 34'b0100111111111010110001000011110011  ;
REGofMAX1DataOut_F4_65 <= 34'b0101000000011110111110110101101001  ;
REGofMAX1DataOut_F4_66 <= 34'b0101000010001001010001101000001111  ;
REGofMAX1DataOut_F4_67 <= 34'b0101000011111010101000101110011110  ;
REGofMAX1DataOut_F4_68 <= 34'b0101000100100010110010111110101110  ;
REGofMAX1DataOut_F4_69 <= 34'b0101000100100001110011110000000000  ;
REGofMAX1DataOut_F4_70 <= 34'b0101000010001010000110100101110110  ;
REGofMAX1DataOut_F4_71 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F4_72 <= 34'b0101000011101110111111001110011011  ;
REGofMAX1DataOut_F4_73 <= 34'b0101000100100000000100001001100111  ;
REGofMAX1DataOut_F4_74 <= 34'b0101000100100010001101010010011010  ;
REGofMAX1DataOut_F4_75 <= 34'b0101000011001101000011011100010001  ;
REGofMAX1DataOut_F4_76 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F4_77 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_78 <= 34'b0100111001011001000100111110011001  ;
REGofMAX1DataOut_F4_79 <= 34'b0101000011100001010010100001011011  ;
REGofMAX1DataOut_F4_80 <= 34'b0101000100011110011101010101100110  ;
REGofMAX1DataOut_F4_81 <= 34'b0101000100100011010110001111001110  ;
REGofMAX1DataOut_F4_82 <= 34'b0101000010100010010010111101010011  ;
REGofMAX1DataOut_F4_83 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F4_84 <= 34'b0101000011100110011101101101101000  ;
REGofMAX1DataOut_F4_85 <= 34'b0101000100011111001011010110001000  ;
REGofMAX1DataOut_F4_86 <= 34'b0101000100100011111101101101100011  ;
REGofMAX1DataOut_F4_87 <= 34'b0101000100000111011010000111001111  ;
REGofMAX1DataOut_F4_88 <= 34'b0101000001010011000111011101010111  ;
REGofMAX1DataOut_F4_89 <= 34'b0101000001100001000101100001100100  ;
REGofMAX1DataOut_F4_90 <= 34'b0101000011001010101001011001111100  ;
REGofMAX1DataOut_F4_91 <= 34'b0101000100000110100111101010111110  ;
REGofMAX1DataOut_F4_92 <= 34'b0101000100011111001001001111001000  ;
REGofMAX1DataOut_F4_93 <= 34'b0101000100011010110000111010011100  ;
REGofMAX1DataOut_F4_94 <= 34'b0101000001011000001101110000110011  ;
REGofMAX1DataOut_F4_95 <= 34'b0000000000000000000000000000000000  ;
REGofMAX1DataOut_F4_96 <= 34'b0101000010110010111011000111000101  ;
REGofMAX1DataOut_F4_97 <= 34'b0101000100000110100001001100111100  ;
REGofMAX1DataOut_F4_98 <= 34'b0101000100011110110101100001001000  ;
REGofMAX1DataOut_F4_99 <= 34'b0101000100011100110010111010110101  ;
REGofMAX1DataOut_F4_100 <= 34'b0101000100000100001010100000000101 ;
REGofMAX1DataOut_F4_101 <= 34'b0101000011110110110110111101100000 ;
REGofMAX1DataOut_F4_102 <= 34'b0101000100000011110111110100100100 ;
REGofMAX1DataOut_F4_103 <= 34'b0101000100010100011011101000100111 ;
REGofMAX1DataOut_F4_104 <= 34'b0101000100011011100010010101111110 ;
REGofMAX1DataOut_F4_105 <= 34'b0101000011111000111111101001001011 ;
REGofMAX1DataOut_F4_106 <= 34'b0000000000000000000000000000000000 ;
REGofMAX1DataOut_F4_107 <= 34'b0100111111101110000010110011011101 ;
REGofMAX1DataOut_F4_108 <= 34'b0101000000100110101100101000000001 ;
REGofMAX1DataOut_F4_109 <= 34'b0101000011011010100001111011011110 ; 
REGofMAX1DataOut_F4_110 <= 34'b0101000100010100011001000000100110 ; 
REGofMAX1DataOut_F4_111 <= 34'b0101000100100000100110010101101110 ; 
REGofMAX1DataOut_F4_112 <= 34'b0101000100011001100101111010110011 ; 
REGofMAX1DataOut_F4_113 <= 34'b0101000100010010000011111101010010 ; 
REGofMAX1DataOut_F4_114 <= 34'b0101000100001011001111110101101100 ; 
REGofMAX1DataOut_F4_115 <= 34'b0101000100001111011100010111001111 ; 
REGofMAX1DataOut_F4_116 <= 34'b0101000100000100100000010001010001 ; 
REGofMAX1DataOut_F4_117 <= 34'b0101000001111110100101110010011101 ; 
REGofMAX1DataOut_F4_118 <= 34'b0000000000000000000000000000000000 ; 
REGofMAX1DataOut_F4_119 <= 34'b0100111111111010010010010001001110 ; 
REGofMAX1DataOut_F4_120 <= 34'b0100111001011001000100111110011001 ;
REGofMAX1DataOut_F4_121 <= 34'b0101000001110111011101101100101010 ; 
REGofMAX1DataOut_F4_122 <= 34'b0101000011100110101110110101110110 ; 
REGofMAX1DataOut_F4_123 <= 34'b0101000100001010111000111101101001 ; 
REGofMAX1DataOut_F4_124 <= 34'b0101000100001111000101111001010111 ; 
REGofMAX1DataOut_F4_125 <= 34'b0101000100001010110111010010011101 ; 
REGofMAX1DataOut_F4_126 <= 34'b0101000100000010111110110100001110 ; 
REGofMAX1DataOut_F4_127 <= 34'b0101000011110000001110100100000000 ; 
REGofMAX1DataOut_F4_128 <= 34'b0101000011001101111100011011000011 ; 
REGofMAX1DataOut_F4_129 <= 34'b0101000001101100100010000111001101 ; 
REGofMAX1DataOut_F4_130 <= 34'b0101000001010011111011011000101110 ; 
REGofMAX1DataOut_F4_131 <= 34'b0100111001011001000100111110011001 ; 
REGofMAX1DataOut_F4_132 <= 34'b0100111001011001000100111110011001 ; 
REGofMAX1DataOut_F4_133 <= 34'b0100111001011001000100111110011001 ; 
REGofMAX1DataOut_F4_134 <= 34'b0101000010011111110011010010110010 ; 
REGofMAX1DataOut_F4_135 <= 34'b0101000011010101110011101001011110 ; 
REGofMAX1DataOut_F4_136 <= 34'b0101000011110000101111101010011001 ; 
REGofMAX1DataOut_F4_137 <= 34'b0101000011110011111000011100010010 ; 
REGofMAX1DataOut_F4_138 <= 34'b0101000011101000011111000001110101 ; 
REGofMAX1DataOut_F4_139 <= 34'b0101000011010111010100001100101110 ; 
REGofMAX1DataOut_F4_140 <= 34'b0101000010101101010011001101010101 ; 
REGofMAX1DataOut_F4_141 <= 34'b0101000001110011110011111100111100 ; 
REGofMAX1DataOut_F4_142 <= 34'b0100111001011001000100111110011001 ; 
REGofMAX1DataOut_F4_143 <= 34'b0100111001011001000100111110011001 ; 


#period;
end 
endmodule




//module 


module happyTB();
reg clk, Conv2LayerStart, inputAXIstart,rst_Controller ;



reg [31:0] AXIinput;
wire [31:0] AXIoutput;

localparam period = 100; 

 
 //happy  happyInstance (clk, rst_Controller, Conv2LayerStart,  AXIinput, AXIoutput, inputAXIstart  );
 happy  happyInstance (clk,  AXIinput, AXIoutput  );
 
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	
//Conv2LayerStart <= 1'b0;
//rst_Controller <= 1'b0;
//inputAXIstart  <= 1'b1;



AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000010001001001010011000 ;
#100;
AXIinput  <=  32'b10010001010000110110101011101110 ;
#100;
AXIinput  <=  32'b10101011010100001110110101110001 ;
#100;
AXIinput  <=  32'b10100110010101000011110111111001 ;
#100;
AXIinput  <=  32'b10111001110001010000111110111111 ;
#100;
AXIinput  <=  32'b10111101111101010100001110010011 ;
#100;
AXIinput  <=  32'b00110010101001000101000010100001 ;
#100;
AXIinput  <=  32'b11010001111101010101010000000110 ;
#100;
AXIinput  <=  32'b00100011010010011010000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000010100 ;
#100;
AXIinput  <=  32'b00100000100101001010111111000101 ;
#100;
AXIinput  <=  32'b00001110010001100011001110101101 ;
#100;
AXIinput  <=  32'b01000100000000001110000111010010 ;
#100;
AXIinput  <=  32'b01010001000001011001001001011110 ;
#100;
AXIinput  <=  32'b11010100010000101000111100001111 ;
#100;
AXIinput  <=  32'b11100101000100001100010110010100 ;
#100;
AXIinput  <=  32'b10101101010001000011000011101011 ;
#100;
AXIinput  <=  32'b11000110010100010000010011001011 ;
#100;
AXIinput  <=  32'b10010111110101000011001011110101 ;
#100;
AXIinput  <=  32'b10000000000101010000010111110011 ;
#100;
AXIinput  <=  32'b00001000100011000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001010000110100 ;
#100;
AXIinput  <=  32'b11001111111100000010010100001110 ;
#100;
AXIinput  <=  32'b01101000000000000110000101000011 ;
#100;
AXIinput  <=  32'b11010001010101101111111101010000 ;
#100;
AXIinput  <=  32'b11110101110000101000011001010100 ;
#100;
AXIinput  <=  32'b00110101000010011111111011010101 ;
#100;
AXIinput  <=  32'b00001110111110010011001111001001 ;
#100;
AXIinput  <=  32'b01000100000111100100011110100010 ;
#100;
AXIinput  <=  32'b01010001000010011101010010010000 ;
#100;
AXIinput  <=  32'b10010100001111111110001111010010 ;
#100;
AXIinput  <=  32'b10010101000011001010110010011101 ;
#100;
AXIinput  <=  32'b01010000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000010100000110100000100000 ;
#100;
AXIinput  <=  32'b00010110010101000011010000100000 ;
#100;
AXIinput  <=  32'b11110100000001010000110110110011 ;
#100;
AXIinput  <=  32'b11100111100010010100001011011010 ;
#100;
AXIinput  <=  32'b01111101000001110000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000101000001 ;
#100;
AXIinput  <=  32'b01011111111101110101110101010000 ;
#100;
AXIinput  <=  32'b11111101011000011111011100010100 ;
#100;
AXIinput  <=  32'b00111111111011100100101010000101 ;
#100;
AXIinput  <=  32'b00001110100111000010100110011101 ;
#100;
AXIinput  <=  32'b01000010000101101110111111110100 ;
#100;
AXIinput  <=  32'b01010000100011010001110110010011 ;
#100;
AXIinput  <=  32'b10010100001100000100110100010010 ;
#100;
AXIinput  <=  32'b11110101000011001000001000110010 ;
#100;
AXIinput  <=  32'b10011101010000101011101101101010 ;
#100;
AXIinput  <=  32'b11110110010100000101000011110100 ;
#100;
AXIinput  <=  32'b10100101000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001010000001111001111 ;
#100;
AXIinput  <=  32'b11110101000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000101000010110010 ;
#100;
AXIinput  <=  32'b10001111000011100001010000111011 ;
#100;
AXIinput  <=  32'b11011110111111000011010100001110 ;
#100;
AXIinput  <=  32'b11011000110000011110000101000010 ;
#100;
AXIinput  <=  32'b11011101111001101110111001010000 ;
#100;
AXIinput  <=  32'b10111111010010110011100101010100 ;
#100;
AXIinput  <=  32'b00110001111001110111001011100101 ;
#100;
AXIinput  <=  32'b00001100110011010001010000111101 ;
#100;
AXIinput  <=  32'b01000011011000110010001100011100 ;
#100;
AXIinput  <=  32'b01010000110011001101110011111111 ;
#100;
AXIinput  <=  32'b10010100000011111111000101000101 ;
#100;
AXIinput  <=  32'b01010000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000101000011100010100111 ;
#100;
AXIinput  <=  32'b10011011110001010000111001110010 ;
#100;
AXIinput  <=  32'b00001101000010010100001100111010 ;
#100;
AXIinput  <=  32'b10010111111000000101000010100010 ;
#100;
AXIinput  <=  32'b10101100001111111101010000110001 ;
#100;
AXIinput  <=  32'b01101010000100010101010100001110 ;
#100;
AXIinput  <=  32'b00110010111111000011100101000011 ;
#100;
AXIinput  <=  32'b10100001011101101001111101010000 ;
#100;
AXIinput  <=  32'b11010100010010000110011111010011 ;
#100;
AXIinput  <=  32'b11111001111100011100001000110000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b01000010011001011000110111000110 ;
#100;
AXIinput  <=  32'b01010000100101100111110001101011 ;
#100;
AXIinput  <=  32'b00010100001100011100001110001110 ;
#100;
AXIinput  <=  32'b00110101000011100010010111011101 ;
#100;
AXIinput  <=  32'b01011001010000110011111000111001 ;
#100;
AXIinput  <=  32'b11001111000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001010000111001001010 ;
#100;
AXIinput  <=  32'b11110011010010010100010000010000 ;
#100;
AXIinput  <=  32'b00111110000011100101000100000010 ;
#100;
AXIinput  <=  32'b00110011000000111001010000110010 ;
#100;
AXIinput  <=  32'b11010011101101001011010100001100 ;
#100;
AXIinput  <=  32'b00001101110011011001010101000011 ;
#100;
AXIinput  <=  32'b10010101111110100011001101010000 ;
#100;
AXIinput  <=  32'b11100010101110100011011001010100 ;
#100;
AXIinput  <=  32'b00101000111100011110001000100101 ;
#100;
AXIinput  <=  32'b00001100011010111010011100001101 ;
#100;
AXIinput  <=  32'b01000011000010001011110000110010 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000001010001000000101111000011 ;
#100;
AXIinput  <=  32'b00001101010100010000101100001011 ;
#100;
AXIinput  <=  32'b00100100110101000100001100011101 ;
#100;
AXIinput  <=  32'b11010111011001010001000010010100 ;
#100;
AXIinput  <=  32'b01101100111000010100010000001110 ;
#100;
AXIinput  <=  32'b00110101001010110101000011110001 ;
#100;
AXIinput  <=  32'b11010110011001000001010000101100 ;
#100;
AXIinput  <=  32'b00000100000101101011010100001010 ;
#100;
AXIinput  <=  32'b00111101011011111010100101000010 ;
#100;
AXIinput  <=  32'b00000001111001010000011000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b01000010100101101101011111101010 ;
#100;
AXIinput  <=  32'b01010001000000100000100000100001 ;
#100;
AXIinput  <=  32'b10010100010000101110000100101011 ;
#100;
AXIinput  <=  32'b01000101000100001011001100100110 ;
#100;
AXIinput  <=  32'b01000001010001000000011111001011 ;
#100;
AXIinput  <=  32'b00101000010100001011000101101000 ;
#100;
AXIinput  <=  32'b10001010000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001010000100100001001 ;
#100;
AXIinput  <=  32'b11010000010100010100000001100111 ;
#100;
AXIinput  <=  32'b10000010110111110000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00010100000100110110110001111110 ;
#100;
AXIinput  <=  32'b00110101000001010100100001101010 ;
#100;
AXIinput  <=  32'b10001100000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000101000000 ;
#100;
AXIinput  <=  32'b00010010010100100000011001010000 ;
#100;
AXIinput  <=  32'b01001000111111101110011010010100 ;
#100;
AXIinput  <=  32'b00011001101010000101101011110000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000001101001000011101000 ;
#100;
AXIinput  <=  32'b01110001010000110011011100001110 ;
#100;
AXIinput  <=  32'b10110100010100001110100001110111 ;
#100;
AXIinput  <=  32'b00000010000101000011101101001110 ;
#100;
AXIinput  <=  32'b10011100100001010000111010111110 ;
#100;
AXIinput  <=  32'b10011111111000010100001110000010 ;
#100;
AXIinput  <=  32'b11011100010011110101000010011111 ;
#100;
AXIinput  <=  32'b10001000001111101001001111001101 ;
#100;
AXIinput  <=  32'b00100000011101011111000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000010100 ;
#100;
AXIinput  <=  32'b00010010111110101111101000100101 ;
#100;
AXIinput  <=  32'b00001011101010110100010110111101 ;
#100;
AXIinput  <=  32'b01000011100010011000001101000001 ;
#100;
AXIinput  <=  32'b01010000110111011000010001111100 ;
#100;
AXIinput  <=  32'b10010100001100010111101000010110 ;
#100;
AXIinput  <=  32'b01100101000011100101011000000011 ;
#100;
AXIinput  <=  32'b10000001010000111011100000010011 ;
#100;
AXIinput  <=  32'b11010100010100001110110111101100 ;
#100;
AXIinput  <=  32'b01001111110101000011000101100100 ;
#100;
AXIinput  <=  32'b11001010010001001111111010111011 ;
#100;
AXIinput  <=  32'b11100010011100000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001010000100111 ;
#100;
AXIinput  <=  32'b11110011110000000101010100000110 ;
#100;
AXIinput  <=  32'b11110100111000011001110000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b01010000111010010111110001110010 ;
#100;
AXIinput  <=  32'b00010100001110010010110100101010 ;
#100;
AXIinput  <=  32'b10000101000010110100011110111111 ;
#100;
AXIinput  <=  32'b01100000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000010100000100000010010101 ;
#100;
AXIinput  <=  32'b11101001110000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001010000101111 ;
#100;
AXIinput  <=  32'b01011000100100001110010100001100 ;
#100;
AXIinput  <=  32'b00011011000100100111000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000010100 ;
#100;
AXIinput  <=  32'b00110100010101100101110111110101 ;
#100;
AXIinput  <=  32'b00001100111101010110010001110001 ;
#100;
AXIinput  <=  32'b01000000110011001100000101001111 ;
#100;
AXIinput  <=  32'b01010000010000100111101110010110 ;
#100;
AXIinput  <=  32'b10000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000010100110011101000111 ;
#100;
AXIinput  <=  32'b10011101010000110101000000101011 ;
#100;
AXIinput  <=  32'b11101110010100001100111110000011 ;
#100;
AXIinput  <=  32'b10001111010101000010101101011001 ;
#100;
AXIinput  <=  32'b00011001010001010000110101000010 ;
#100;
AXIinput  <=  32'b01011101011111010100001011101110 ;
#100;
AXIinput  <=  32'b10101110001010000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001010000100000 ;
#100;
AXIinput  <=  32'b10100101110110000001010100001011 ;
#100;
AXIinput  <=  32'b10011100000010010000100101000010 ;
#100;
AXIinput  <=  32'b00100111101111111010111101010000 ;
#100;
AXIinput  <=  32'b01011110101011000000100010010100 ;
#100;
AXIinput  <=  32'b00101011010000111001111010110101 ;
#100;
AXIinput  <=  32'b00001010110000110100011011111001 ;
#100;
AXIinput  <=  32'b01000010101011111101011110101000 ;
#100;
AXIinput  <=  32'b01010000100010110101001110000100 ;
#100;
AXIinput  <=  32'b01000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000010100010100101101000 ;
#100;
AXIinput  <=  32'b10100001010000110011000110010110 ;
#100;
AXIinput  <=  32'b11101000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001010000101101100111 ;
#100;
AXIinput  <=  32'b01110010110000010100001001000001 ;
#100;
AXIinput  <=  32'b00001010000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000010100000110 ;
#100;
AXIinput  <=  32'b10101100110010110010110101000010 ;
#100;
AXIinput  <=  32'b11010110100110111100000101010000 ;
#100;
AXIinput  <=  32'b10110100111111000010100110000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b01000010110000111000111101001011 ;
#100;
AXIinput  <=  32'b01010000101110111000011101000011 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000010010101010010010000 ;
#100;
AXIinput  <=  32'b00001001010000100101000111011010 ;
#100;
AXIinput  <=  32'b00110101010100001010100101010100 ;
#100;
AXIinput  <=  32'b01101101100000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000010100001101011110 ;
#100;
AXIinput  <=  32'b10000101011010000101000011100110 ;
#100;
AXIinput  <=  32'b01010000110011011001010000110000 ;
#100;
AXIinput  <=  32'b01111011000011010011010100001010 ;
#100;
AXIinput  <=  32'b01111111101101001011100101000011 ;
#100;
AXIinput  <=  32'b00001010101001110110111101010000 ;
#100;
AXIinput  <=  32'b11001101111011010101010000010100 ;
#100;
AXIinput  <=  32'b00100010101111100101011110110000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b01000001100110010001111000001000 ;
#100;
AXIinput  <=  32'b01010000101001010100100000001000 ;
#100;
AXIinput  <=  32'b00010100001100000000111110000110 ;
#100;
AXIinput  <=  32'b01000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000010100001110111000001001 ;
#100;
AXIinput  <=  32'b01111010000101000011110001011010 ;
#100;
AXIinput  <=  32'b10000100001101010000111010010101 ;
#100;
AXIinput  <=  32'b11011111011001010100001101100011 ;
#100;
AXIinput  <=  32'b11101101110100100101000010010000 ;
#100;
AXIinput  <=  32'b10100110011001111001010000100111 ;
#100;
AXIinput  <=  32'b10010111111110010001010011111110 ;
#100;
AXIinput  <=  32'b10100011110000100111000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000001010000 ;
#100;
AXIinput  <=  32'b01000000010100100001101101010100 ;
#100;
AXIinput  <=  32'b00110001100010101010110001010101 ;
#100;
AXIinput  <=  32'b00001100001100110101101011011000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001010000100011 ;
#100;
AXIinput  <=  32'b10011101111100011010010100001100 ;
#100;
AXIinput  <=  32'b10100000101011010011110101000011 ;
#100;
AXIinput  <=  32'b00010011001001000000111000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b01000001110001010010111001100001 ;
#100;
AXIinput  <=  32'b01010000100011111001000111001101 ;
#100;
AXIinput  <=  32'b10010100000110101111100100101011 ;
#100;
AXIinput  <=  32'b10100000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001010000101100111111 ;
#100;
AXIinput  <=  32'b01110100101000010100001110000111 ;
#100;
AXIinput  <=  32'b00000011111110000101000011100101 ;
#100;
AXIinput  <=  32'b01010100101001100001010000111001 ;
#100;
AXIinput  <=  32'b11101101100010000001010100001101 ;
#100;
AXIinput  <=  32'b01110010111000010100100101000011 ;
#100;
AXIinput  <=  32'b00111110101100010000001001010000 ;
#100;
AXIinput  <=  32'b10011010001110100110001101000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b01001110110011101100010111001110 ;
#100;
AXIinput  <=  32'b01010011101100111011000101110011 ;
#100;
AXIinput  <=  32'b10010101000010000010011111001100 ;
#100;
AXIinput  <=  32'b00011001010000110011110110010001 ;
#100;
AXIinput  <=  32'b11010101010100001110011101100011 ;
#100;
AXIinput  <=  32'b01011110010101000011101100011011 ;
#100;
AXIinput  <=  32'b00010000101101010000111010011110 ;
#100;
AXIinput  <=  32'b00101111100011010100001100010001 ;
#100;
AXIinput  <=  32'b01001111100001000101000000001110 ;
#100;
AXIinput  <=  32'b00100100010101100101001110110011 ;
#100;
AXIinput  <=  32'b10110001011100111001010011101100 ;
#100;
AXIinput  <=  32'b11101100010111001110010100111011 ;
#100;
AXIinput  <=  32'b00111011000101110011100101001110 ;
#100;
AXIinput  <=  32'b11001110110001011100111001010100 ;
#100;
AXIinput  <=  32'b00011111001111110001101111110101 ;
#100;
AXIinput  <=  32'b00001110110001010110010001101101 ;
#100;
AXIinput  <=  32'b01000100000011111111010100010110 ;
#100;
AXIinput  <=  32'b01010001000100011101111110110111 ;
#100;
AXIinput  <=  32'b11010100010001111001111100000000 ;
#100;
AXIinput  <=  32'b10110101000100100010111011010010 ;
#100;
AXIinput  <=  32'b00100101010001001000001110001001 ;
#100;
AXIinput  <=  32'b11101011010100010000001111100110 ;
#100;
AXIinput  <=  32'b10110011110101000010101001111111 ;
#100;
AXIinput  <=  32'b00100101010101001110110011101100 ;
#100;
AXIinput  <=  32'b01011100111001010011101100111011 ;
#100;
AXIinput  <=  32'b00010111001110010100111011001110 ;
#100;
AXIinput  <=  32'b11000101110011100101010000110110 ;
#100;
AXIinput  <=  32'b11101011101110001100010100001111 ;
#100;
AXIinput  <=  32'b01010001010101101001000101000100 ;
#100;
AXIinput  <=  32'b00110101001111001001110101010001 ;
#100;
AXIinput  <=  32'b00100001101010101110100011010100 ;
#100;
AXIinput  <=  32'b01001001000000100001010101010101 ;
#100;
AXIinput  <=  32'b00010010101001110001101010010001 ;
#100;
AXIinput  <=  32'b01000100101101110001100001000000 ;
#100;
AXIinput  <=  32'b01010001001011011001110000011111 ;
#100;
AXIinput  <=  32'b10010100010000111101000001000001 ;
#100;
AXIinput  <=  32'b10010101000010111011011111011011 ;
#100;
AXIinput  <=  32'b10100001001110110011101100010111 ;
#100;
AXIinput  <=  32'b00111001010100000110001000010101 ;
#100;
AXIinput  <=  32'b01001000100101000011100111000101 ;
#100;
AXIinput  <=  32'b01101010100101010000111101001110 ;
#100;
AXIinput  <=  32'b10000011000110010100010001001011 ;
#100;
AXIinput  <=  32'b11000000110010110101000100011101 ;
#100;
AXIinput  <=  32'b10001001000101000101010001000101 ;
#100;
AXIinput  <=  32'b00010100110010001011010100010000 ;
#100;
AXIinput  <=  32'b11000010101110100000110101000100 ;
#100;
AXIinput  <=  32'b10010111010100111010000101010001 ;
#100;
AXIinput  <=  32'b00101101001101100010111110010100 ;
#100;
AXIinput  <=  32'b01001010111000100110000110010101 ;
#100;
AXIinput  <=  32'b00010000010010010010010001001101 ;
#100;
AXIinput  <=  32'b00111011001110110001011100111001 ;
#100;
AXIinput  <=  32'b01010000100110001111010101100000 ;
#100;
AXIinput  <=  32'b10010100001101110011001100010011 ;
#100;
AXIinput  <=  32'b01010101000100001001100101000110 ;
#100;
AXIinput  <=  32'b11111001010001000110010110001111 ;
#100;
AXIinput  <=  32'b00110100010100010000011101000100 ;
#100;
AXIinput  <=  32'b01001100100101000011111011010011 ;
#100;
AXIinput  <=  32'b11011000111001010000110000111011 ;
#100;
AXIinput  <=  32'b01111111110000010100001110100111 ;
#100;
AXIinput  <=  32'b10110010100101110101000100100100 ;
#100;
AXIinput  <=  32'b11111111100110110101010001001010 ;
#100;
AXIinput  <=  32'b11100100100111011111010100010001 ;
#100;
AXIinput  <=  32'b11000100011100110110110101000010 ;
#100;
AXIinput  <=  32'b11111010110000000000101001010000 ;
#100;
AXIinput  <=  32'b11000100010011000001001000010100 ;
#100;
AXIinput  <=  32'b00111000011100100001010111100101 ;
#100;
AXIinput  <=  32'b00010001110011101001010001110101 ;
#100;
AXIinput  <=  32'b01000100100011010111011110111011 ;
#100;
AXIinput  <=  32'b01010000111110001101101010001101 ;
#100;
AXIinput  <=  32'b01010100000110110011111110000101 ;
#100;
AXIinput  <=  32'b01010100111011001110110001011100 ;
#100;
AXIinput  <=  32'b11100100000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000010100010000010111100111 ;
#100;
AXIinput  <=  32'b00100000000101000100101000001010 ;
#100;
AXIinput  <=  32'b11100100000101010001001000101110 ;
#100;
AXIinput  <=  32'b00011011011001010100001110010000 ;
#100;
AXIinput  <=  32'b01100010001110100101000011000100 ;
#100;
AXIinput  <=  32'b11111000000100111101010000111011 ;
#100;
AXIinput  <=  32'b00110010011100001111010100010010 ;
#100;
AXIinput  <=  32'b01110000110000101101110101000100 ;
#100;
AXIinput  <=  32'b10010111100100000111010101010000 ;
#100;
AXIinput  <=  32'b11110110000011100000000111010011 ;
#100;
AXIinput  <=  32'b10110011101100010111001110010100 ;
#100;
AXIinput  <=  32'b11101100111011000101110011100101 ;
#100;
AXIinput  <=  32'b01000001110100111110110101000011 ;
#100;
AXIinput  <=  32'b01010000111000000011010001001110 ;
#100;
AXIinput  <=  32'b01010100010010001011010010110111 ;
#100;
AXIinput  <=  32'b11100101000100100011101110111000 ;
#100;
AXIinput  <=  32'b11100101010000111101001110110000 ;
#100;
AXIinput  <=  32'b00110111000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000101000011100110100100 ;
#100;
AXIinput  <=  32'b01011001011001010001001010010100 ;
#100;
AXIinput  <=  32'b10010111001001010100010010111010 ;
#100;
AXIinput  <=  32'b00111000101100000101000100010001 ;
#100;
AXIinput  <=  32'b10010001011100001001010000101010 ;
#100;
AXIinput  <=  32'b10110110011100000011010100001010 ;
#100;
AXIinput  <=  32'b11111010110011101101000101000011 ;
#100;
AXIinput  <=  32'b10101111111101011011101101010000 ;
#100;
AXIinput  <=  32'b11101001000000001000100101010100 ;
#100;
AXIinput  <=  32'b01000100110100110100111101100101 ;
#100;
AXIinput  <=  32'b00010010001001011010001010101001 ;
#100;
AXIinput  <=  32'b01000011110100111011000010100001 ;
#100;
AXIinput  <=  32'b01001110110011101100010111001110 ;
#100;
AXIinput  <=  32'b01000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000100011110000101011101 ;
#100;
AXIinput  <=  32'b11110101010001001011101000010101 ;
#100;
AXIinput  <=  32'b00010011010100010010110111011011 ;
#100;
AXIinput  <=  32'b10000101100101000100011100000101 ;
#100;
AXIinput  <=  32'b01110011100001010001000001111100 ;
#100;
AXIinput  <=  32'b00101100100110010100010000010011 ;
#100;
AXIinput  <=  32'b00101100001101100101000100001000 ;
#100;
AXIinput  <=  32'b01001111101110110101010001000111 ;
#100;
AXIinput  <=  32'b10100010101101101001010100010001 ;
#100;
AXIinput  <=  32'b10100000101110100000000101000011 ;
#100;
AXIinput  <=  32'b01001111101001011010111101001110 ;
#100;
AXIinput  <=  32'b11001110110001011100111001000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000101 ;
#100;
AXIinput  <=  32'b00001101110001001001010001000101 ;
#100;
AXIinput  <=  32'b01000100100101000110100111101100 ;
#100;
AXIinput  <=  32'b01010001001011101010100100011101 ;
#100;
AXIinput  <=  32'b10010100010010101101100000010100 ;
#100;
AXIinput  <=  32'b11000101000100100100101011111011 ;
#100;
AXIinput  <=  32'b10001001010001000110011100100101 ;
#100;
AXIinput  <=  32'b10010010010100010001011111001110 ;
#100;
AXIinput  <=  32'b11011001000101000100011011101011 ;
#100;
AXIinput  <=  32'b11101001101001010001000010100100 ;
#100;
AXIinput  <=  32'b00010001001110010100000100100110 ;
#100;
AXIinput  <=  32'b10010000011000100100111011001110 ;
#100;
AXIinput  <=  32'b11000101110011100101001110110011 ;
#100;
AXIinput  <=  32'b10110001011100111001000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000101000011 ;
#100;
AXIinput  <=  32'b01111001000101001001111101010001 ;
#100;
AXIinput  <=  32'b00011100001010110010110010010100 ;
#100;
AXIinput  <=  32'b01001000101000111010001101000101 ;
#100;
AXIinput  <=  32'b00010010001000011000010110000101 ;
#100;
AXIinput  <=  32'b01000100011000001110101010001010 ;
#100;
AXIinput  <=  32'b01010001000100100000110011001100 ;
#100;
AXIinput  <=  32'b01010100010000101111111110010011 ;
#100;
AXIinput  <=  32'b11100101000011010001000110010000 ;
#100;
AXIinput  <=  32'b11100001001110110011101100010111 ;
#100;
AXIinput  <=  32'b00111001010011101100111011000101 ;
#100;
AXIinput  <=  32'b11001110010100111011001110110001 ;
#100;
AXIinput  <=  32'b01110011100101001110110011101100 ;
#100;
AXIinput  <=  32'b01011100111001000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000101000010001001 ;
#100;
AXIinput  <=  32'b10110101010001111001010000111001 ;
#100;
AXIinput  <=  32'b01101001101011101011010100001111 ;
#100;
AXIinput  <=  32'b10101111101111111010000101000011 ;
#100;
AXIinput  <=  32'b11101010100010100100000101010000 ;
#100;
AXIinput  <=  32'b11101001010001000000011110010100 ;
#100;
AXIinput  <=  32'b00110000001000111011110010000100 ;
#100;
AXIinput  <=  32'b11101100111011000101110011100101 ;
#100;
AXIinput  <=  32'b00111011001110110001011100111001 ;
#100;
AXIinput  <=  32'b01001110010110010001001111100110 ;
#100;
AXIinput  <=  32'b01010011100101100100010011111001 ;
#100;
AXIinput  <=  32'b10010101000010011011001001100000 ;
#100;
AXIinput  <=  32'b10101001010000111001101001011001 ;
#100;
AXIinput  <=  32'b00111000010100001111101000010011 ;
#100;
AXIinput  <=  32'b00001111000101000011111110010001 ;
#100;
AXIinput  <=  32'b11000001011001010000111011001111 ;
#100;
AXIinput  <=  32'b11011011000111010100001010100001 ;
#100;
AXIinput  <=  32'b10110000111110000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001001110010110 ;
#100;
AXIinput  <=  32'b01000100111110011001010011100101 ;
#100;
AXIinput  <=  32'b10010001001111100110010100111001 ;
#100;
AXIinput  <=  32'b01100100010011111001100101001110 ;
#100;
AXIinput  <=  32'b01011001000100111110011001010100 ;
#100;
AXIinput  <=  32'b00100101010001001100000111110101 ;
#100;
AXIinput  <=  32'b00010000000000001010001111001101 ;
#100;
AXIinput  <=  32'b01000100010000011101000001010001 ;
#100;
AXIinput  <=  32'b01010001000011110001000110001101 ;
#100;
AXIinput  <=  32'b11010100010000110001100000010100 ;
#100;
AXIinput  <=  32'b01110101000100000111011101011110 ;
#100;
AXIinput  <=  32'b10101001010000111101111000101000 ;
#100;
AXIinput  <=  32'b01110000010100001011100010111101 ;
#100;
AXIinput  <=  32'b00111111000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001001110010110010001 ;
#100;
AXIinput  <=  32'b00111110011001010011100101100100 ;
#100;
AXIinput  <=  32'b01001111100110010100111001011001 ;
#100;
AXIinput  <=  32'b00010011111001100101010000111100 ;
#100;
AXIinput  <=  32'b00000000111010010010010100010001 ;
#100;
AXIinput  <=  32'b10001110101101100000100101000100 ;
#100;
AXIinput  <=  32'b01110101001101100110010001010001 ;
#100;
AXIinput  <=  32'b00010101000101111111100001010100 ;
#100;
AXIinput  <=  32'b01000010100000100010001100100101 ;
#100;
AXIinput  <=  32'b00010000111111010000101010101001 ;
#100;
AXIinput  <=  32'b01000100010100011000110000001111 ;
#100;
AXIinput  <=  32'b01010001000001100101110000010011 ;
#100;
AXIinput  <=  32'b01000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000001001110010110010001001111 ;
#100;
AXIinput  <=  32'b10011001010100000111101101111010 ;
#100;
AXIinput  <=  32'b10111101000101000100001100101111 ;
#100;
AXIinput  <=  32'b01001011111101010001000111010001 ;
#100;
AXIinput  <=  32'b00101111000000010100010001001001 ;
#100;
AXIinput  <=  32'b00111001001011010101000100000000 ;
#100;
AXIinput  <=  32'b01100111111001111001010000111010 ;
#100;
AXIinput  <=  32'b01110000000001100111010100010000 ;
#100;
AXIinput  <=  32'b10101001010001001011100101000100 ;
#100;
AXIinput  <=  32'b01110110100100101001010001010001 ;
#100;
AXIinput  <=  32'b00011111101011011100110110010100 ;
#100;
AXIinput  <=  32'b00111101010110100100011000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b00111001011001000100111110011001 ;
#100;
AXIinput  <=  32'b01010000101100001001010011100100 ;
#100;
AXIinput  <=  32'b01010100010001100000000110001111 ;
#100;
AXIinput  <=  32'b11000101000100100000101111111100 ;
#100;
AXIinput  <=  32'b10110101010000111011010111100100 ;
#100;
AXIinput  <=  32'b10101000010100001100010101110000 ;
#100;
AXIinput  <=  32'b11011101100101000011000101110000 ;
#100;
AXIinput  <=  32'b00101110110001010000111001010001 ;
#100;
AXIinput  <=  32'b10010100110010010100010001011101 ;
#100;
AXIinput  <=  32'b11001010111100000101000100100010 ;
#100;
AXIinput  <=  32'b00001010001100100101010001000100 ;
#100;
AXIinput  <=  32'b10111101100111111011000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000100111001 ;
#100;
AXIinput  <=  32'b01100100010011111001100101010000 ;
#100;
AXIinput  <=  32'b11101101100101101111101010010100 ;
#100;
AXIinput  <=  32'b01000111110111110001010011010101 ;
#100;
AXIinput  <=  32'b00010010001010111001010001111001 ;
#100;
AXIinput  <=  32'b01000010110111101101100000010000 ;
#100;
AXIinput  <=  32'b01001111111110101100010000111100 ;
#100;
AXIinput  <=  32'b11010100000001111011111011010110 ;
#100;
AXIinput  <=  32'b10010101000010001001010001101000 ;
#100;
AXIinput  <=  32'b00111101010000111110101010001011 ;
#100;
AXIinput  <=  32'b10011110010100010010001011001011 ;
#100;
AXIinput  <=  32'b11101011100101000100100001110011 ;
#100;
AXIinput  <=  32'b11000000000001010000100010100001 ;
#100;
AXIinput  <=  32'b10100101110110000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000101000011101110 ;
#100;
AXIinput  <=  32'b11111100111001101101010001001000 ;
#100;
AXIinput  <=  32'b00000100001001100111010100010010 ;
#100;
AXIinput  <=  32'b00100011010100100110100101000011 ;
#100;
AXIinput  <=  32'b00110100001101110001000100000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000010011 ;
#100;
AXIinput  <=  32'b10010110010001001111100110010100 ;
#100;
AXIinput  <=  32'b11100101100100010011111001100101 ;
#100;
AXIinput  <=  32'b01000011100001010010100001011011 ;
#100;
AXIinput  <=  32'b01010001000111100111010101011001 ;
#100;
AXIinput  <=  32'b10010100010010001101011000111100 ;
#100;
AXIinput  <=  32'b11100101000010100010010010111101 ;
#100;
AXIinput  <=  32'b01001100000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000010100001110011001110110 ;
#100;
AXIinput  <=  32'b11011010000101000100011111001011 ;
#100;
AXIinput  <=  32'b01011000100001010001001000111111 ;
#100;
AXIinput  <=  32'b01101101100011010100010000011101 ;
#100;
AXIinput  <=  32'b10100001110011110101000001010011 ;
#100;
AXIinput  <=  32'b00011101110101011101010000011000 ;
#100;
AXIinput  <=  32'b01000101100001100100010100001100 ;
#100;
AXIinput  <=  32'b10101010010110011111000101000100 ;
#100;
AXIinput  <=  32'b00011010011110101011111001010001 ;
#100;
AXIinput  <=  32'b00011111001001001111001000010100 ;
#100;
AXIinput  <=  32'b01000110101100001110100111000101 ;
#100;
AXIinput  <=  32'b00000101100000110111000011001100 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b01010000101100101110110001110001 ;
#100;
AXIinput  <=  32'b01010100010000011010000100110011 ;
#100;
AXIinput  <=  32'b11000101000100011110110101100001 ;
#100;
AXIinput  <=  32'b00100001010001000111001100101110 ;
#100;
AXIinput  <=  32'b10110101010100010000010000101010 ;
#100;
AXIinput  <=  32'b00000001010101000011110110110110 ;
#100;
AXIinput  <=  32'b11110110000001010001000000111101 ;
#100;
AXIinput  <=  32'b11110100100100010100010001010001 ;
#100;
AXIinput  <=  32'b10111010001001110101000100011011 ;
#100;
AXIinput  <=  32'b10001001010111111001010000111110 ;
#100;
AXIinput  <=  32'b00111111101001001011000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000100111111 ;
#100;
AXIinput  <=  32'b10111000001011001101110101010000 ;
#100;
AXIinput  <=  32'b00100110101100101000000001010100 ;
#100;
AXIinput  <=  32'b00110110101000011110110111100101 ;
#100;
AXIinput  <=  32'b00010001010001100100000010011001 ;
#100;
AXIinput  <=  32'b01000100100000100110010101101110 ;
#100;
AXIinput  <=  32'b01010001000110011001011110101100 ;
#100;
AXIinput  <=  32'b11010100010001001000001111110101 ;
#100;
AXIinput  <=  32'b00100101000100001011001111110101 ;
#100;
AXIinput  <=  32'b10110001010001000011110111000101 ;
#100;
AXIinput  <=  32'b11001111010100010000010010000001 ;
#100;
AXIinput  <=  32'b00010100010101000001111110100101 ;
#100;
AXIinput  <=  32'b11001001110100000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000010011111111101001 ;
#100;
AXIinput  <=  32'b00100100010011100100111001011001 ;
#100;
AXIinput  <=  32'b00010011111001100101010000011101 ;
#100;
AXIinput  <=  32'b11011101101100101010010100001110 ;
#100;
AXIinput  <=  32'b01101011101101011101100101000100 ;
#100;
AXIinput  <=  32'b00101011100011110110100101010001 ;
#100;
AXIinput  <=  32'b00001111000101111001010111010100 ;
#100;
AXIinput  <=  32'b01000010101101110100100111010101 ;
#100;
AXIinput  <=  32'b00010000001011111011010000111001 ;
#100;
AXIinput  <=  32'b01000011110000001110100100000000 ;
#100;
AXIinput  <=  32'b01010000110011011111000110110000 ;
#100;
AXIinput  <=  32'b11010100000110110010001000011100 ;
#100;
AXIinput  <=  32'b11010101000001010011111011011000 ;
#100;
AXIinput  <=  32'b10111001001110010110010001001111 ;
#100;
AXIinput  <=  32'b10011001010011100101100100010011 ;
#100;
AXIinput  <=  32'b11100110010100111001011001000100 ;
#100;
AXIinput  <=  32'b11111001100101010000100111111100 ;
#100;
AXIinput  <=  32'b11010010110010010100001101010111 ;
#100;
AXIinput  <=  32'b00111010010111100101000011110000 ;
#100;
AXIinput  <=  32'b10111110101001100101010000111100 ;
#100;
AXIinput  <=  32'b11111000011100010010010100001110 ;
#100;
AXIinput  <=  32'b10000111110000011101010101000011 ;
#100;
AXIinput  <=  32'b01011101010000110010111001010000 ;
#100;
AXIinput  <=  32'b10101101010011001101010101010100 ;
#100;
AXIinput  <=  32'b00011100111100111111001111000100 ;
#100;
AXIinput  <=  32'b11100101100100010011111001100101 ;
#100;
AXIinput  <=  32'b00111001011001000100111110011001 ;
#100;

//Conv2LayerStart <= 1'b1;
//inputAXIstart <= 1'b0;
 

#period;
end 
endmodule






module AXIinputhappyTB();
reg clk, AXIstart, Conv2LayerStart ; 
wire MAX2LayerFinish;
reg [31:0] AXIinput;

wire [33:0] REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143 ;

wire [33:0] MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 ;

localparam period = 100; 

 
 AXIinputFromARM_3_1  AXIinstance (clk, AXIinput, AXIstart , 
REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143 
);

MERGEHOPE_L3_L4 l3_l4instance (clk, Conv2LayerStart, MAX2LayerFinish
,REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143 
,MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 
 );
 
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	
AXIstart <= 1'b1;
Conv2LayerStart <= 1'b0;


AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000010001001001010011000 ;
#100;
AXIinput  <=  32'b10010001010000110110101011101110 ;
#100;
AXIinput  <=  32'b10101011010100001110110101110001 ;
#100;
AXIinput  <=  32'b10100110010101000011110111111001 ;
#100;
AXIinput  <=  32'b10111001110001010000111110111111 ;
#100;
AXIinput  <=  32'b10111101111101010100001110010011 ;
#100;
AXIinput  <=  32'b00110010101001000101000010100001 ;
#100;
AXIinput  <=  32'b11010001111101010101010000000110 ;
#100;
AXIinput  <=  32'b00100011010010011010000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000010100 ;
#100;
AXIinput  <=  32'b00100000100101001010111111000101 ;
#100;
AXIinput  <=  32'b00001110010001100011001110101101 ;
#100;
AXIinput  <=  32'b01000100000000001110000111010010 ;
#100;
AXIinput  <=  32'b01010001000001011001001001011110 ;
#100;
AXIinput  <=  32'b11010100010000101000111100001111 ;
#100;
AXIinput  <=  32'b11100101000100001100010110010100 ;
#100;
AXIinput  <=  32'b10101101010001000011000011101011 ;
#100;
AXIinput  <=  32'b11000110010100010000010011001011 ;
#100;
AXIinput  <=  32'b10010111110101000011001011110101 ;
#100;
AXIinput  <=  32'b10000000000101010000010111110011 ;
#100;
AXIinput  <=  32'b00001000100011000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001010000110100 ;
#100;
AXIinput  <=  32'b11001111111100000010010100001110 ;
#100;
AXIinput  <=  32'b01101000000000000110000101000011 ;
#100;
AXIinput  <=  32'b11010001010101101111111101010000 ;
#100;
AXIinput  <=  32'b11110101110000101000011001010100 ;
#100;
AXIinput  <=  32'b00110101000010011111111011010101 ;
#100;
AXIinput  <=  32'b00001110111110010011001111001001 ;
#100;
AXIinput  <=  32'b01000100000111100100011110100010 ;
#100;
AXIinput  <=  32'b01010001000010011101010010010000 ;
#100;
AXIinput  <=  32'b10010100001111111110001111010010 ;
#100;
AXIinput  <=  32'b10010101000011001010110010011101 ;
#100;
AXIinput  <=  32'b01010000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000010100000110100000100000 ;
#100;
AXIinput  <=  32'b00010110010101000011010000100000 ;
#100;
AXIinput  <=  32'b11110100000001010000110110110011 ;
#100;
AXIinput  <=  32'b11100111100010010100001011011010 ;
#100;
AXIinput  <=  32'b01111101000001110000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000101000001 ;
#100;
AXIinput  <=  32'b01011111111101110101110101010000 ;
#100;
AXIinput  <=  32'b11111101011000011111011100010100 ;
#100;
AXIinput  <=  32'b00111111111011100100101010000101 ;
#100;
AXIinput  <=  32'b00001110100111000010100110011101 ;
#100;
AXIinput  <=  32'b01000010000101101110111111110100 ;
#100;
AXIinput  <=  32'b01010000100011010001110110010011 ;
#100;
AXIinput  <=  32'b10010100001100000100110100010010 ;
#100;
AXIinput  <=  32'b11110101000011001000001000110010 ;
#100;
AXIinput  <=  32'b10011101010000101011101101101010 ;
#100;
AXIinput  <=  32'b11110110010100000101000011110100 ;
#100;
AXIinput  <=  32'b10100101000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001010000001111001111 ;
#100;
AXIinput  <=  32'b11110101000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000101000010110010 ;
#100;
AXIinput  <=  32'b10001111000011100001010000111011 ;
#100;
AXIinput  <=  32'b11011110111111000011010100001110 ;
#100;
AXIinput  <=  32'b11011000110000011110000101000010 ;
#100;
AXIinput  <=  32'b11011101111001101110111001010000 ;
#100;
AXIinput  <=  32'b10111111010010110011100101010100 ;
#100;
AXIinput  <=  32'b00110001111001110111001011100101 ;
#100;
AXIinput  <=  32'b00001100110011010001010000111101 ;
#100;
AXIinput  <=  32'b01000011011000110010001100011100 ;
#100;
AXIinput  <=  32'b01010000110011001101110011111111 ;
#100;
AXIinput  <=  32'b10010100000011111111000101000101 ;
#100;
AXIinput  <=  32'b01010000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000101000011100010100111 ;
#100;
AXIinput  <=  32'b10011011110001010000111001110010 ;
#100;
AXIinput  <=  32'b00001101000010010100001100111010 ;
#100;
AXIinput  <=  32'b10010111111000000101000010100010 ;
#100;
AXIinput  <=  32'b10101100001111111101010000110001 ;
#100;
AXIinput  <=  32'b01101010000100010101010100001110 ;
#100;
AXIinput  <=  32'b00110010111111000011100101000011 ;
#100;
AXIinput  <=  32'b10100001011101101001111101010000 ;
#100;
AXIinput  <=  32'b11010100010010000110011111010011 ;
#100;
AXIinput  <=  32'b11111001111100011100001000110000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b01000010011001011000110111000110 ;
#100;
AXIinput  <=  32'b01010000100101100111110001101011 ;
#100;
AXIinput  <=  32'b00010100001100011100001110001110 ;
#100;
AXIinput  <=  32'b00110101000011100010010111011101 ;
#100;
AXIinput  <=  32'b01011001010000110011111000111001 ;
#100;
AXIinput  <=  32'b11001111000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001010000111001001010 ;
#100;
AXIinput  <=  32'b11110011010010010100010000010000 ;
#100;
AXIinput  <=  32'b00111110000011100101000100000010 ;
#100;
AXIinput  <=  32'b00110011000000111001010000110010 ;
#100;
AXIinput  <=  32'b11010011101101001011010100001100 ;
#100;
AXIinput  <=  32'b00001101110011011001010101000011 ;
#100;
AXIinput  <=  32'b10010101111110100011001101010000 ;
#100;
AXIinput  <=  32'b11100010101110100011011001010100 ;
#100;
AXIinput  <=  32'b00101000111100011110001000100101 ;
#100;
AXIinput  <=  32'b00001100011010111010011100001101 ;
#100;
AXIinput  <=  32'b01000011000010001011110000110010 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000001010001000000101111000011 ;
#100;
AXIinput  <=  32'b00001101010100010000101100001011 ;
#100;
AXIinput  <=  32'b00100100110101000100001100011101 ;
#100;
AXIinput  <=  32'b11010111011001010001000010010100 ;
#100;
AXIinput  <=  32'b01101100111000010100010000001110 ;
#100;
AXIinput  <=  32'b00110101001010110101000011110001 ;
#100;
AXIinput  <=  32'b11010110011001000001010000101100 ;
#100;
AXIinput  <=  32'b00000100000101101011010100001010 ;
#100;
AXIinput  <=  32'b00111101011011111010100101000010 ;
#100;
AXIinput  <=  32'b00000001111001010000011000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b01000010100101101101011111101010 ;
#100;
AXIinput  <=  32'b01010001000000100000100000100001 ;
#100;
AXIinput  <=  32'b10010100010000101110000100101011 ;
#100;
AXIinput  <=  32'b01000101000100001011001100100110 ;
#100;
AXIinput  <=  32'b01000001010001000000011111001011 ;
#100;
AXIinput  <=  32'b00101000010100001011000101101000 ;
#100;
AXIinput  <=  32'b10001010000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001010000100100001001 ;
#100;
AXIinput  <=  32'b11010000010100010100000001100111 ;
#100;
AXIinput  <=  32'b10000010110111110000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00010100000100110110110001111110 ;
#100;
AXIinput  <=  32'b00110101000001010100100001101010 ;
#100;
AXIinput  <=  32'b10001100000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000101000000 ;
#100;
AXIinput  <=  32'b00010010010100100000011001010000 ;
#100;
AXIinput  <=  32'b01001000111111101110011010010100 ;
#100;
AXIinput  <=  32'b00011001101010000101101011110000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000001101001000011101000 ;
#100;
AXIinput  <=  32'b01110001010000110011011100001110 ;
#100;
AXIinput  <=  32'b10110100010100001110100001110111 ;
#100;
AXIinput  <=  32'b00000010000101000011101101001110 ;
#100;
AXIinput  <=  32'b10011100100001010000111010111110 ;
#100;
AXIinput  <=  32'b10011111111000010100001110000010 ;
#100;
AXIinput  <=  32'b11011100010011110101000010011111 ;
#100;
AXIinput  <=  32'b10001000001111101001001111001101 ;
#100;
AXIinput  <=  32'b00100000011101011111000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000010100 ;
#100;
AXIinput  <=  32'b00010010111110101111101000100101 ;
#100;
AXIinput  <=  32'b00001011101010110100010110111101 ;
#100;
AXIinput  <=  32'b01000011100010011000001101000001 ;
#100;
AXIinput  <=  32'b01010000110111011000010001111100 ;
#100;
AXIinput  <=  32'b10010100001100010111101000010110 ;
#100;
AXIinput  <=  32'b01100101000011100101011000000011 ;
#100;
AXIinput  <=  32'b10000001010000111011100000010011 ;
#100;
AXIinput  <=  32'b11010100010100001110110111101100 ;
#100;
AXIinput  <=  32'b01001111110101000011000101100100 ;
#100;
AXIinput  <=  32'b11001010010001001111111010111011 ;
#100;
AXIinput  <=  32'b11100010011100000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001010000100111 ;
#100;
AXIinput  <=  32'b11110011110000000101010100000110 ;
#100;
AXIinput  <=  32'b11110100111000011001110000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b01010000111010010111110001110010 ;
#100;
AXIinput  <=  32'b00010100001110010010110100101010 ;
#100;
AXIinput  <=  32'b10000101000010110100011110111111 ;
#100;
AXIinput  <=  32'b01100000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000010100000100000010010101 ;
#100;
AXIinput  <=  32'b11101001110000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001010000101111 ;
#100;
AXIinput  <=  32'b01011000100100001110010100001100 ;
#100;
AXIinput  <=  32'b00011011000100100111000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000010100 ;
#100;
AXIinput  <=  32'b00110100010101100101110111110101 ;
#100;
AXIinput  <=  32'b00001100111101010110010001110001 ;
#100;
AXIinput  <=  32'b01000000110011001100000101001111 ;
#100;
AXIinput  <=  32'b01010000010000100111101110010110 ;
#100;
AXIinput  <=  32'b10000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000010100110011101000111 ;
#100;
AXIinput  <=  32'b10011101010000110101000000101011 ;
#100;
AXIinput  <=  32'b11101110010100001100111110000011 ;
#100;
AXIinput  <=  32'b10001111010101000010101101011001 ;
#100;
AXIinput  <=  32'b00011001010001010000110101000010 ;
#100;
AXIinput  <=  32'b01011101011111010100001011101110 ;
#100;
AXIinput  <=  32'b10101110001010000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001010000100000 ;
#100;
AXIinput  <=  32'b10100101110110000001010100001011 ;
#100;
AXIinput  <=  32'b10011100000010010000100101000010 ;
#100;
AXIinput  <=  32'b00100111101111111010111101010000 ;
#100;
AXIinput  <=  32'b01011110101011000000100010010100 ;
#100;
AXIinput  <=  32'b00101011010000111001111010110101 ;
#100;
AXIinput  <=  32'b00001010110000110100011011111001 ;
#100;
AXIinput  <=  32'b01000010101011111101011110101000 ;
#100;
AXIinput  <=  32'b01010000100010110101001110000100 ;
#100;
AXIinput  <=  32'b01000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000010100010100101101000 ;
#100;
AXIinput  <=  32'b10100001010000110011000110010110 ;
#100;
AXIinput  <=  32'b11101000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001010000101101100111 ;
#100;
AXIinput  <=  32'b01110010110000010100001001000001 ;
#100;
AXIinput  <=  32'b00001010000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000010100000110 ;
#100;
AXIinput  <=  32'b10101100110010110010110101000010 ;
#100;
AXIinput  <=  32'b11010110100110111100000101010000 ;
#100;
AXIinput  <=  32'b10110100111111000010100110000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b01000010110000111000111101001011 ;
#100;
AXIinput  <=  32'b01010000101110111000011101000011 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000010010101010010010000 ;
#100;
AXIinput  <=  32'b00001001010000100101000111011010 ;
#100;
AXIinput  <=  32'b00110101010100001010100101010100 ;
#100;
AXIinput  <=  32'b01101101100000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000010100001101011110 ;
#100;
AXIinput  <=  32'b10000101011010000101000011100110 ;
#100;
AXIinput  <=  32'b01010000110011011001010000110000 ;
#100;
AXIinput  <=  32'b01111011000011010011010100001010 ;
#100;
AXIinput  <=  32'b01111111101101001011100101000011 ;
#100;
AXIinput  <=  32'b00001010101001110110111101010000 ;
#100;
AXIinput  <=  32'b11001101111011010101010000010100 ;
#100;
AXIinput  <=  32'b00100010101111100101011110110000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b01000001100110010001111000001000 ;
#100;
AXIinput  <=  32'b01010000101001010100100000001000 ;
#100;
AXIinput  <=  32'b00010100001100000000111110000110 ;
#100;
AXIinput  <=  32'b01000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000010100001110111000001001 ;
#100;
AXIinput  <=  32'b01111010000101000011110001011010 ;
#100;
AXIinput  <=  32'b10000100001101010000111010010101 ;
#100;
AXIinput  <=  32'b11011111011001010100001101100011 ;
#100;
AXIinput  <=  32'b11101101110100100101000010010000 ;
#100;
AXIinput  <=  32'b10100110011001111001010000100111 ;
#100;
AXIinput  <=  32'b10010111111110010001010011111110 ;
#100;
AXIinput  <=  32'b10100011110000100111000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000001010000 ;
#100;
AXIinput  <=  32'b01000000010100100001101101010100 ;
#100;
AXIinput  <=  32'b00110001100010101010110001010101 ;
#100;
AXIinput  <=  32'b00001100001100110101101011011000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001010000100011 ;
#100;
AXIinput  <=  32'b10011101111100011010010100001100 ;
#100;
AXIinput  <=  32'b10100000101011010011110101000011 ;
#100;
AXIinput  <=  32'b00010011001001000000111000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b01000001110001010010111001100001 ;
#100;
AXIinput  <=  32'b01010000100011111001000111001101 ;
#100;
AXIinput  <=  32'b10010100000110101111100100101011 ;
#100;
AXIinput  <=  32'b10100000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001010000101100111111 ;
#100;
AXIinput  <=  32'b01110100101000010100001110000111 ;
#100;
AXIinput  <=  32'b00000011111110000101000011100101 ;
#100;
AXIinput  <=  32'b01010100101001100001010000111001 ;
#100;
AXIinput  <=  32'b11101101100010000001010100001101 ;
#100;
AXIinput  <=  32'b01110010111000010100100101000011 ;
#100;
AXIinput  <=  32'b00111110101100010000001001010000 ;
#100;
AXIinput  <=  32'b10011010001110100110001101000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b01001110110011101100010111001110 ;
#100;
AXIinput  <=  32'b01010011101100111011000101110011 ;
#100;
AXIinput  <=  32'b10010101000010000010011111001100 ;
#100;
AXIinput  <=  32'b00011001010000110011110110010001 ;
#100;
AXIinput  <=  32'b11010101010100001110011101100011 ;
#100;
AXIinput  <=  32'b01011110010101000011101100011011 ;
#100;
AXIinput  <=  32'b00010000101101010000111010011110 ;
#100;
AXIinput  <=  32'b00101111100011010100001100010001 ;
#100;
AXIinput  <=  32'b01001111100001000101000000001110 ;
#100;
AXIinput  <=  32'b00100100010101100101001110110011 ;
#100;
AXIinput  <=  32'b10110001011100111001010011101100 ;
#100;
AXIinput  <=  32'b11101100010111001110010100111011 ;
#100;
AXIinput  <=  32'b00111011000101110011100101001110 ;
#100;
AXIinput  <=  32'b11001110110001011100111001010100 ;
#100;
AXIinput  <=  32'b00011111001111110001101111110101 ;
#100;
AXIinput  <=  32'b00001110110001010110010001101101 ;
#100;
AXIinput  <=  32'b01000100000011111111010100010110 ;
#100;
AXIinput  <=  32'b01010001000100011101111110110111 ;
#100;
AXIinput  <=  32'b11010100010001111001111100000000 ;
#100;
AXIinput  <=  32'b10110101000100100010111011010010 ;
#100;
AXIinput  <=  32'b00100101010001001000001110001001 ;
#100;
AXIinput  <=  32'b11101011010100010000001111100110 ;
#100;
AXIinput  <=  32'b10110011110101000010101001111111 ;
#100;
AXIinput  <=  32'b00100101010101001110110011101100 ;
#100;
AXIinput  <=  32'b01011100111001010011101100111011 ;
#100;
AXIinput  <=  32'b00010111001110010100111011001110 ;
#100;
AXIinput  <=  32'b11000101110011100101010000110110 ;
#100;
AXIinput  <=  32'b11101011101110001100010100001111 ;
#100;
AXIinput  <=  32'b01010001010101101001000101000100 ;
#100;
AXIinput  <=  32'b00110101001111001001110101010001 ;
#100;
AXIinput  <=  32'b00100001101010101110100011010100 ;
#100;
AXIinput  <=  32'b01001001000000100001010101010101 ;
#100;
AXIinput  <=  32'b00010010101001110001101010010001 ;
#100;
AXIinput  <=  32'b01000100101101110001100001000000 ;
#100;
AXIinput  <=  32'b01010001001011011001110000011111 ;
#100;
AXIinput  <=  32'b10010100010000111101000001000001 ;
#100;
AXIinput  <=  32'b10010101000010111011011111011011 ;
#100;
AXIinput  <=  32'b10100001001110110011101100010111 ;
#100;
AXIinput  <=  32'b00111001010100000110001000010101 ;
#100;
AXIinput  <=  32'b01001000100101000011100111000101 ;
#100;
AXIinput  <=  32'b01101010100101010000111101001110 ;
#100;
AXIinput  <=  32'b10000011000110010100010001001011 ;
#100;
AXIinput  <=  32'b11000000110010110101000100011101 ;
#100;
AXIinput  <=  32'b10001001000101000101010001000101 ;
#100;
AXIinput  <=  32'b00010100110010001011010100010000 ;
#100;
AXIinput  <=  32'b11000010101110100000110101000100 ;
#100;
AXIinput  <=  32'b10010111010100111010000101010001 ;
#100;
AXIinput  <=  32'b00101101001101100010111110010100 ;
#100;
AXIinput  <=  32'b01001010111000100110000110010101 ;
#100;
AXIinput  <=  32'b00010000010010010010010001001101 ;
#100;
AXIinput  <=  32'b00111011001110110001011100111001 ;
#100;
AXIinput  <=  32'b01010000100110001111010101100000 ;
#100;
AXIinput  <=  32'b10010100001101110011001100010011 ;
#100;
AXIinput  <=  32'b01010101000100001001100101000110 ;
#100;
AXIinput  <=  32'b11111001010001000110010110001111 ;
#100;
AXIinput  <=  32'b00110100010100010000011101000100 ;
#100;
AXIinput  <=  32'b01001100100101000011111011010011 ;
#100;
AXIinput  <=  32'b11011000111001010000110000111011 ;
#100;
AXIinput  <=  32'b01111111110000010100001110100111 ;
#100;
AXIinput  <=  32'b10110010100101110101000100100100 ;
#100;
AXIinput  <=  32'b11111111100110110101010001001010 ;
#100;
AXIinput  <=  32'b11100100100111011111010100010001 ;
#100;
AXIinput  <=  32'b11000100011100110110110101000010 ;
#100;
AXIinput  <=  32'b11111010110000000000101001010000 ;
#100;
AXIinput  <=  32'b11000100010011000001001000010100 ;
#100;
AXIinput  <=  32'b00111000011100100001010111100101 ;
#100;
AXIinput  <=  32'b00010001110011101001010001110101 ;
#100;
AXIinput  <=  32'b01000100100011010111011110111011 ;
#100;
AXIinput  <=  32'b01010000111110001101101010001101 ;
#100;
AXIinput  <=  32'b01010100000110110011111110000101 ;
#100;
AXIinput  <=  32'b01010100111011001110110001011100 ;
#100;
AXIinput  <=  32'b11100100000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000010100010000010111100111 ;
#100;
AXIinput  <=  32'b00100000000101000100101000001010 ;
#100;
AXIinput  <=  32'b11100100000101010001001000101110 ;
#100;
AXIinput  <=  32'b00011011011001010100001110010000 ;
#100;
AXIinput  <=  32'b01100010001110100101000011000100 ;
#100;
AXIinput  <=  32'b11111000000100111101010000111011 ;
#100;
AXIinput  <=  32'b00110010011100001111010100010010 ;
#100;
AXIinput  <=  32'b01110000110000101101110101000100 ;
#100;
AXIinput  <=  32'b10010111100100000111010101010000 ;
#100;
AXIinput  <=  32'b11110110000011100000000111010011 ;
#100;
AXIinput  <=  32'b10110011101100010111001110010100 ;
#100;
AXIinput  <=  32'b11101100111011000101110011100101 ;
#100;
AXIinput  <=  32'b01000001110100111110110101000011 ;
#100;
AXIinput  <=  32'b01010000111000000011010001001110 ;
#100;
AXIinput  <=  32'b01010100010010001011010010110111 ;
#100;
AXIinput  <=  32'b11100101000100100011101110111000 ;
#100;
AXIinput  <=  32'b11100101010000111101001110110000 ;
#100;
AXIinput  <=  32'b00110111000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000101000011100110100100 ;
#100;
AXIinput  <=  32'b01011001011001010001001010010100 ;
#100;
AXIinput  <=  32'b10010111001001010100010010111010 ;
#100;
AXIinput  <=  32'b00111000101100000101000100010001 ;
#100;
AXIinput  <=  32'b10010001011100001001010000101010 ;
#100;
AXIinput  <=  32'b10110110011100000011010100001010 ;
#100;
AXIinput  <=  32'b11111010110011101101000101000011 ;
#100;
AXIinput  <=  32'b10101111111101011011101101010000 ;
#100;
AXIinput  <=  32'b11101001000000001000100101010100 ;
#100;
AXIinput  <=  32'b01000100110100110100111101100101 ;
#100;
AXIinput  <=  32'b00010010001001011010001010101001 ;
#100;
AXIinput  <=  32'b01000011110100111011000010100001 ;
#100;
AXIinput  <=  32'b01001110110011101100010111001110 ;
#100;
AXIinput  <=  32'b01000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000101000100011110000101011101 ;
#100;
AXIinput  <=  32'b11110101010001001011101000010101 ;
#100;
AXIinput  <=  32'b00010011010100010010110111011011 ;
#100;
AXIinput  <=  32'b10000101100101000100011100000101 ;
#100;
AXIinput  <=  32'b01110011100001010001000001111100 ;
#100;
AXIinput  <=  32'b00101100100110010100010000010011 ;
#100;
AXIinput  <=  32'b00101100001101100101000100001000 ;
#100;
AXIinput  <=  32'b01001111101110110101010001000111 ;
#100;
AXIinput  <=  32'b10100010101101101001010100010001 ;
#100;
AXIinput  <=  32'b10100000101110100000000101000011 ;
#100;
AXIinput  <=  32'b01001111101001011010111101001110 ;
#100;
AXIinput  <=  32'b11001110110001011100111001000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000101 ;
#100;
AXIinput  <=  32'b00001101110001001001010001000101 ;
#100;
AXIinput  <=  32'b01000100100101000110100111101100 ;
#100;
AXIinput  <=  32'b01010001001011101010100100011101 ;
#100;
AXIinput  <=  32'b10010100010010101101100000010100 ;
#100;
AXIinput  <=  32'b11000101000100100100101011111011 ;
#100;
AXIinput  <=  32'b10001001010001000110011100100101 ;
#100;
AXIinput  <=  32'b10010010010100010001011111001110 ;
#100;
AXIinput  <=  32'b11011001000101000100011011101011 ;
#100;
AXIinput  <=  32'b11101001101001010001000010100100 ;
#100;
AXIinput  <=  32'b00010001001110010100000100100110 ;
#100;
AXIinput  <=  32'b10010000011000100100111011001110 ;
#100;
AXIinput  <=  32'b11000101110011100101001110110011 ;
#100;
AXIinput  <=  32'b10110001011100111001000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000101000011 ;
#100;
AXIinput  <=  32'b01111001000101001001111101010001 ;
#100;
AXIinput  <=  32'b00011100001010110010110010010100 ;
#100;
AXIinput  <=  32'b01001000101000111010001101000101 ;
#100;
AXIinput  <=  32'b00010010001000011000010110000101 ;
#100;
AXIinput  <=  32'b01000100011000001110101010001010 ;
#100;
AXIinput  <=  32'b01010001000100100000110011001100 ;
#100;
AXIinput  <=  32'b01010100010000101111111110010011 ;
#100;
AXIinput  <=  32'b11100101000011010001000110010000 ;
#100;
AXIinput  <=  32'b11100001001110110011101100010111 ;
#100;
AXIinput  <=  32'b00111001010011101100111011000101 ;
#100;
AXIinput  <=  32'b11001110010100111011001110110001 ;
#100;
AXIinput  <=  32'b01110011100101001110110011101100 ;
#100;
AXIinput  <=  32'b01011100111001000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000101000010001001 ;
#100;
AXIinput  <=  32'b10110101010001111001010000111001 ;
#100;
AXIinput  <=  32'b01101001101011101011010100001111 ;
#100;
AXIinput  <=  32'b10101111101111111010000101000011 ;
#100;
AXIinput  <=  32'b11101010100010100100000101010000 ;
#100;
AXIinput  <=  32'b11101001010001000000011110010100 ;
#100;
AXIinput  <=  32'b00110000001000111011110010000100 ;
#100;
AXIinput  <=  32'b11101100111011000101110011100101 ;
#100;
AXIinput  <=  32'b00111011001110110001011100111001 ;
#100;
AXIinput  <=  32'b01001110010110010001001111100110 ;
#100;
AXIinput  <=  32'b01010011100101100100010011111001 ;
#100;
AXIinput  <=  32'b10010101000010011011001001100000 ;
#100;
AXIinput  <=  32'b10101001010000111001101001011001 ;
#100;
AXIinput  <=  32'b00111000010100001111101000010011 ;
#100;
AXIinput  <=  32'b00001111000101000011111110010001 ;
#100;
AXIinput  <=  32'b11000001011001010000111011001111 ;
#100;
AXIinput  <=  32'b11011011000111010100001010100001 ;
#100;
AXIinput  <=  32'b10110000111110000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000001001110010110 ;
#100;
AXIinput  <=  32'b01000100111110011001010011100101 ;
#100;
AXIinput  <=  32'b10010001001111100110010100111001 ;
#100;
AXIinput  <=  32'b01100100010011111001100101001110 ;
#100;
AXIinput  <=  32'b01011001000100111110011001010100 ;
#100;
AXIinput  <=  32'b00100101010001001100000111110101 ;
#100;
AXIinput  <=  32'b00010000000000001010001111001101 ;
#100;
AXIinput  <=  32'b01000100010000011101000001010001 ;
#100;
AXIinput  <=  32'b01010001000011110001000110001101 ;
#100;
AXIinput  <=  32'b11010100010000110001100000010100 ;
#100;
AXIinput  <=  32'b01110101000100000111011101011110 ;
#100;
AXIinput  <=  32'b10101001010000111101111000101000 ;
#100;
AXIinput  <=  32'b01110000010100001011100010111101 ;
#100;
AXIinput  <=  32'b00111111000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000001001110010110010001 ;
#100;
AXIinput  <=  32'b00111110011001010011100101100100 ;
#100;
AXIinput  <=  32'b01001111100110010100111001011001 ;
#100;
AXIinput  <=  32'b00010011111001100101010000111100 ;
#100;
AXIinput  <=  32'b00000000111010010010010100010001 ;
#100;
AXIinput  <=  32'b10001110101101100000100101000100 ;
#100;
AXIinput  <=  32'b01110101001101100110010001010001 ;
#100;
AXIinput  <=  32'b00010101000101111111100001010100 ;
#100;
AXIinput  <=  32'b01000010100000100010001100100101 ;
#100;
AXIinput  <=  32'b00010000111111010000101010101001 ;
#100;
AXIinput  <=  32'b01000100010100011000110000001111 ;
#100;
AXIinput  <=  32'b01010001000001100101110000010011 ;
#100;
AXIinput  <=  32'b01000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000001001110010110010001001111 ;
#100;
AXIinput  <=  32'b10011001010100000111101101111010 ;
#100;
AXIinput  <=  32'b10111101000101000100001100101111 ;
#100;
AXIinput  <=  32'b01001011111101010001000111010001 ;
#100;
AXIinput  <=  32'b00101111000000010100010001001001 ;
#100;
AXIinput  <=  32'b00111001001011010101000100000000 ;
#100;
AXIinput  <=  32'b01100111111001111001010000111010 ;
#100;
AXIinput  <=  32'b01110000000001100111010100010000 ;
#100;
AXIinput  <=  32'b10101001010001001011100101000100 ;
#100;
AXIinput  <=  32'b01110110100100101001010001010001 ;
#100;
AXIinput  <=  32'b00011111101011011100110110010100 ;
#100;
AXIinput  <=  32'b00111101010110100100011000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000001 ;
#100;
AXIinput  <=  32'b00111001011001000100111110011001 ;
#100;
AXIinput  <=  32'b01010000101100001001010011100100 ;
#100;
AXIinput  <=  32'b01010100010001100000000110001111 ;
#100;
AXIinput  <=  32'b11000101000100100000101111111100 ;
#100;
AXIinput  <=  32'b10110101010000111011010111100100 ;
#100;
AXIinput  <=  32'b10101000010100001100010101110000 ;
#100;
AXIinput  <=  32'b11011101100101000011000101110000 ;
#100;
AXIinput  <=  32'b00101110110001010000111001010001 ;
#100;
AXIinput  <=  32'b10010100110010010100010001011101 ;
#100;
AXIinput  <=  32'b11001010111100000101000100100010 ;
#100;
AXIinput  <=  32'b00001010001100100101010001000100 ;
#100;
AXIinput  <=  32'b10111101100111111011000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000100111001 ;
#100;
AXIinput  <=  32'b01100100010011111001100101010000 ;
#100;
AXIinput  <=  32'b11101101100101101111101010010100 ;
#100;
AXIinput  <=  32'b01000111110111110001010011010101 ;
#100;
AXIinput  <=  32'b00010010001010111001010001111001 ;
#100;
AXIinput  <=  32'b01000010110111101101100000010000 ;
#100;
AXIinput  <=  32'b01001111111110101100010000111100 ;
#100;
AXIinput  <=  32'b11010100000001111011111011010110 ;
#100;
AXIinput  <=  32'b10010101000010001001010001101000 ;
#100;
AXIinput  <=  32'b00111101010000111110101010001011 ;
#100;
AXIinput  <=  32'b10011110010100010010001011001011 ;
#100;
AXIinput  <=  32'b11101011100101000100100001110011 ;
#100;
AXIinput  <=  32'b11000000000001010000100010100001 ;
#100;
AXIinput  <=  32'b10100101110110000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000101000011101110 ;
#100;
AXIinput  <=  32'b11111100111001101101010001001000 ;
#100;
AXIinput  <=  32'b00000100001001100111010100010010 ;
#100;
AXIinput  <=  32'b00100011010100100110100101000011 ;
#100;
AXIinput  <=  32'b00110100001101110001000100000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000000010011 ;
#100;
AXIinput  <=  32'b10010110010001001111100110010100 ;
#100;
AXIinput  <=  32'b11100101100100010011111001100101 ;
#100;
AXIinput  <=  32'b01000011100001010010100001011011 ;
#100;
AXIinput  <=  32'b01010001000111100111010101011001 ;
#100;
AXIinput  <=  32'b10010100010010001101011000111100 ;
#100;
AXIinput  <=  32'b11100101000010100010010010111101 ;
#100;
AXIinput  <=  32'b01001100000000000000000000000000 ;
#100;
AXIinput  <=  32'b00000000010100001110011001110110 ;
#100;
AXIinput  <=  32'b11011010000101000100011111001011 ;
#100;
AXIinput  <=  32'b01011000100001010001001000111111 ;
#100;
AXIinput  <=  32'b01101101100011010100010000011101 ;
#100;
AXIinput  <=  32'b10100001110011110101000001010011 ;
#100;
AXIinput  <=  32'b00011101110101011101010000011000 ;
#100;
AXIinput  <=  32'b01000101100001100100010100001100 ;
#100;
AXIinput  <=  32'b10101010010110011111000101000100 ;
#100;
AXIinput  <=  32'b00011010011110101011111001010001 ;
#100;
AXIinput  <=  32'b00011111001001001111001000010100 ;
#100;
AXIinput  <=  32'b01000110101100001110100111000101 ;
#100;
AXIinput  <=  32'b00000101100000110111000011001100 ;
#100;
AXIinput  <=  32'b00000000000000000000000000000000 ;
#100;
AXIinput  <=  32'b01010000101100101110110001110001 ;
#100;
AXIinput  <=  32'b01010100010000011010000100110011 ;
#100;
AXIinput  <=  32'b11000101000100011110110101100001 ;
#100;
AXIinput  <=  32'b00100001010001000111001100101110 ;
#100;
AXIinput  <=  32'b10110101010100010000010000101010 ;
#100;
AXIinput  <=  32'b00000001010101000011110110110110 ;
#100;
AXIinput  <=  32'b11110110000001010001000000111101 ;
#100;
AXIinput  <=  32'b11110100100100010100010001010001 ;
#100;
AXIinput  <=  32'b10111010001001110101000100011011 ;
#100;
AXIinput  <=  32'b10001001010111111001010000111110 ;
#100;
AXIinput  <=  32'b00111111101001001011000000000000 ;
#100;
AXIinput  <=  32'b00000000000000000000000100111111 ;
#100;
AXIinput  <=  32'b10111000001011001101110101010000 ;
#100;
AXIinput  <=  32'b00100110101100101000000001010100 ;
#100;
AXIinput  <=  32'b00110110101000011110110111100101 ;
#100;
AXIinput  <=  32'b00010001010001100100000010011001 ;
#100;
AXIinput  <=  32'b01000100100000100110010101101110 ;
#100;
AXIinput  <=  32'b01010001000110011001011110101100 ;
#100;
AXIinput  <=  32'b11010100010001001000001111110101 ;
#100;
AXIinput  <=  32'b00100101000100001011001111110101 ;
#100;
AXIinput  <=  32'b10110001010001000011110111000101 ;
#100;
AXIinput  <=  32'b11001111010100010000010010000001 ;
#100;
AXIinput  <=  32'b00010100010101000001111110100101 ;
#100;
AXIinput  <=  32'b11001001110100000000000000000000 ;
#100;
AXIinput  <=  32'b00000000000000010011111111101001 ;
#100;
AXIinput  <=  32'b00100100010011100100111001011001 ;
#100;
AXIinput  <=  32'b00010011111001100101010000011101 ;
#100;
AXIinput  <=  32'b11011101101100101010010100001110 ;
#100;
AXIinput  <=  32'b01101011101101011101100101000100 ;
#100;
AXIinput  <=  32'b00101011100011110110100101010001 ;
#100;
AXIinput  <=  32'b00001111000101111001010111010100 ;
#100;
AXIinput  <=  32'b01000010101101110100100111010101 ;
#100;
AXIinput  <=  32'b00010000001011111011010000111001 ;
#100;
AXIinput  <=  32'b01000011110000001110100100000000 ;
#100;
AXIinput  <=  32'b01010000110011011111000110110000 ;
#100;
AXIinput  <=  32'b11010100000110110010001000011100 ;
#100;
AXIinput  <=  32'b11010101000001010011111011011000 ;
#100;
AXIinput  <=  32'b10111001001110010110010001001111 ;
#100;
AXIinput  <=  32'b10011001010011100101100100010011 ;
#100;
AXIinput  <=  32'b11100110010100111001011001000100 ;
#100;
AXIinput  <=  32'b11111001100101010000100111111100 ;
#100;
AXIinput  <=  32'b11010010110010010100001101010111 ;
#100;
AXIinput  <=  32'b00111010010111100101000011110000 ;
#100;
AXIinput  <=  32'b10111110101001100101010000111100 ;
#100;
AXIinput  <=  32'b11111000011100010010010100001110 ;
#100;
AXIinput  <=  32'b10000111110000011101010101000011 ;
#100;
AXIinput  <=  32'b01011101010000110010111001010000 ;
#100;
AXIinput  <=  32'b10101101010011001101010101010100 ;
#100;
AXIinput  <=  32'b00011100111100111111001111000100 ;
#100;
AXIinput  <=  32'b11100101100100010011111001100101 ;
#100;
AXIinput  <=  32'b00111001011001000100111110011001 ;
#100;

Conv2LayerStart <= 1'b1;
AXIstart <= 1'b0;
#period;
end 
endmodule






module AXIoutputTB();


reg clk, outputAXIstart ;
wire [31:0] AXIoutput;

reg [33:0] MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 ;

localparam period = 100; 

 
 AXIoutputToARM_3_1 outputInstance (clk, AXIoutput, outputAXIstart , 
MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 
);

always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
begin	

outputAXIstart  <= 1'b1;


MAX2Data2_OutF4_0   <=  34'b0101000100010110010001011101111011   ;
MAX2Data2_OutF4_1   <=  34'b0101000100101001010000100001001011   ;
MAX2Data2_OutF4_2   <=  34'b0101000100110101101101001101110000   ;
MAX2Data2_OutF4_3   <=  34'b0101000100101000011100111001011010   ;
MAX2Data2_OutF4_4   <=  34'b0101000011001111110100100011100110   ;
MAX2Data2_OutF4_5   <=  34'b0101000100100001100000010111101110   ;
MAX2Data2_OutF4_6   <=  34'b0101000100110010001110111110010011   ;
MAX2Data2_OutF4_7   <=  34'b0101000101000101101011001100110011   ;
MAX2Data2_OutF4_8   <=  34'b0101000101000110100101101100011111   ;
MAX2Data2_OutF4_9   <=  34'b0101000100010110101011110011110101   ;
MAX2Data2_OutF4_10  <=  34'b0101000100110110001000111010101001   ;
MAX2Data2_OutF4_11  <=  34'b0101000100010100000100111101111010   ;
MAX2Data2_OutF4_12  <=  34'b0101000100100001100000011011110111   ;
MAX2Data2_OutF4_13  <=  34'b0101000101000000100100110001000101   ;
MAX2Data2_OutF4_14  <=  34'b0101000100100000001111011011010010   ;
MAX2Data2_OutF4_15  <=  34'b0101000100111110010110000100100110   ;
MAX2Data2_OutF4_16  <=  34'b0101000100101100001000100000001000   ;
MAX2Data2_OutF4_17  <=  34'b0101000100010001101010000001110110   ;
MAX2Data2_OutF4_18  <=  34'b0101000100101111001101111101110101   ;
MAX2Data2_OutF4_19  <=  34'b0101000100011000111100110101101100   ;
MAX2Data2_OutF4_20  <=  34'b0101000101000001110111100110110011   ;
MAX2Data2_OutF4_21  <=  34'b0101000101000011110011000111001000   ;
MAX2Data2_OutF4_22  <=  34'b0101000101000010001001101100100100   ;
MAX2Data2_OutF4_23  <=  34'b0101000100110101011101010011111010   ;
MAX2Data2_OutF4_24  <=  34'b0101000100100010010000011011110111   ;


#period;
end 
endmodule

module ROM_FPGA_Input(out, addr, clk);
output reg [31:0] out;
input[9:0] addr;
input clk;


reg [31:0] ROM[612:0];

initial begin

ROM[0] <=  32'b00000000000000000000000000000000 ; 
ROM[1] <=  32'b00000000000000000000000000000000 ;
ROM[2] <=  32'b00000101000010001001001010011000 ;
ROM[3] <=  32'b10010001010000110110101011101110 ;
ROM[4] <=  32'b10101011010100001110110101110001 ;
ROM[5] <=  32'b10100110010101000011110111111001 ;
ROM[6] <=  32'b10111001110001010000111110111111 ;
ROM[7] <=  32'b10111101111101010100001110010011 ;
ROM[8] <=  32'b00110010101001000101000010100001 ;
ROM[9] <=  32'b11010001111101010101010000000110 ;
ROM[10] <=  32'b00100011010010011010000000000000 ;
ROM[11] <=  32'b00000000000000000000000000000000 ;
ROM[12] <=  32'b00000000000000000000000000000000 ;
ROM[13] <=  32'b00000000000000000000000000010100 ;
ROM[14] <=  32'b00100000100101001010111111000101 ;
ROM[15] <=  32'b00001110010001100011001110101101 ;
ROM[16] <=  32'b01000100000000001110000111010010 ;
ROM[17] <=  32'b01010001000001011001001001011110 ;
ROM[18] <=  32'b11010100010000101000111100001111 ;
ROM[19] <=  32'b11100101000100001100010110010100 ;
ROM[20] <=  32'b10101101010001000011000011101011 ;
ROM[21] <=  32'b11000110010100010000010011001011 ;
ROM[22] <=  32'b10010111110101000011001011110101 ;
ROM[23] <=  32'b10000000000101010000010111110011 ;
ROM[24] <=  32'b00001000100011000000000000000000 ;
ROM[25] <=  32'b00000000000000000000000000000000 ;
ROM[26] <=  32'b00000000000000000001010000110100 ;
ROM[27] <=  32'b11001111111100000010010100001110 ;
ROM[28] <=  32'b01101000000000000110000101000011 ;
ROM[29] <=  32'b11010001010101101111111101010000 ;
ROM[30] <=  32'b11110101110000101000011001010100 ;
ROM[31] <=  32'b00110101000010011111111011010101 ;
ROM[32] <=  32'b00001110111110010011001111001001 ;
ROM[33] <=  32'b01000100000111100100011110100010 ;
ROM[34] <=  32'b01010001000010011101010010010000 ;
ROM[35] <=  32'b10010100001111111110001111010010 ;
ROM[36] <=  32'b10010101000011001010110010011101 ;
ROM[37] <=  32'b01010000000000000000000000000000 ;
ROM[38] <=  32'b00000000010100000110100000100000 ;
ROM[39] <=  32'b00010110010101000011010000100000 ;
ROM[40] <=  32'b11110100000001010000110110110011 ;
ROM[41] <=  32'b11100111100010010100001011011010 ;
ROM[42] <=  32'b01111101000001110000000000000000 ;
ROM[43] <=  32'b00000000000000000000000000000000 ;
ROM[44] <=  32'b00000000000000000000000000000000 ;
ROM[45] <=  32'b00000000000000000000000101000001 ;
ROM[46] <=  32'b01011111111101110101110101010000 ;
ROM[47] <=  32'b11111101011000011111011100010100 ;
ROM[48] <=  32'b00111111111011100100101010000101 ;
ROM[49] <=  32'b00001110100111000010100110011101 ;
ROM[50] <=  32'b01000010000101101110111111110100 ;
ROM[51] <=  32'b01010000100011010001110110010011 ;
ROM[52] <=  32'b10010100001100000100110100010010 ;
ROM[53] <=  32'b11110101000011001000001000110010 ;
ROM[54] <=  32'b10011101010000101011101101101010 ;
ROM[55] <=  32'b11110110010100000101000011110100 ;
ROM[56] <=  32'b10100101000000000000000000000000 ;
ROM[57] <=  32'b00000000000001010000001111001111 ;
ROM[58] <=  32'b11110101000000000000000000000000 ;
ROM[59] <=  32'b00000000000000000101000010110010 ;
ROM[60] <=  32'b10001111000011100001010000111011 ;
ROM[61] <=  32'b11011110111111000011010100001110 ;
ROM[62] <=  32'b11011000110000011110000101000010 ;
ROM[63] <=  32'b11011101111001101110111001010000 ;
ROM[64] <=  32'b10111111010010110011100101010100 ;
ROM[65] <=  32'b00110001111001110111001011100101 ;
ROM[66] <=  32'b00001100110011010001010000111101 ;
ROM[67] <=  32'b01000011011000110010001100011100 ;
ROM[68] <=  32'b01010000110011001101110011111111 ;
ROM[69] <=  32'b10010100000011111111000101000101 ;
ROM[70] <=  32'b01010000000000000000000000000000 ;
ROM[71] <=  32'b00000000000000000000000000000000 ;
ROM[72] <=  32'b00000000000000000000000000000000 ;
ROM[73] <=  32'b00000000000101000011100010100111 ;
ROM[74] <=  32'b10011011110001010000111001110010 ;
ROM[75] <=  32'b00001101000010010100001100111010 ;
ROM[76] <=  32'b10010111111000000101000010100010 ;
ROM[77] <=  32'b10101100001111111101010000110001 ;
ROM[78] <=  32'b01101010000100010101010100001110 ;
ROM[79] <=  32'b00110010111111000011100101000011 ;
ROM[80] <=  32'b10100001011101101001111101010000 ;
ROM[81] <=  32'b11010100010010000110011111010011 ;
ROM[82] <=  32'b11111001111100011100001000110000 ;
ROM[83] <=  32'b00000000000000000000000000000001 ;
ROM[84] <=  32'b01000010011001011000110111000110 ;
ROM[85] <=  32'b01010000100101100111110001101011 ;
ROM[86] <=  32'b00010100001100011100001110001110 ;
ROM[87] <=  32'b00110101000011100010010111011101 ;
ROM[88] <=  32'b01011001010000110011111000111001 ;
ROM[89] <=  32'b11001111000000000000000000000000 ;
ROM[90] <=  32'b00000000000000000000000000000000 ;
ROM[91] <=  32'b00000000000001010000111001001010 ;
ROM[92] <=  32'b11110011010010010100010000010000 ;
ROM[93] <=  32'b00111110000011100101000100000010 ;
ROM[94] <=  32'b00110011000000111001010000110010 ;
ROM[95] <=  32'b11010011101101001011010100001100 ;
ROM[96] <=  32'b00001101110011011001010101000011 ;
ROM[97] <=  32'b10010101111110100011001101010000 ;
ROM[98] <=  32'b11100010101110100011011001010100 ;
ROM[99] <=  32'b00101000111100011110001000100101 ;
ROM[100] <=  32'b00001100011010111010011100001101 ;
ROM[101] <=  32'b01000011000010001011110000110010 ;
ROM[102] <=  32'b00000000000000000000000000000000 ;
ROM[103] <=  32'b00000000000000000000000000000000 ;
ROM[104] <=  32'b00000000000000000000000000000000 ;
ROM[105] <=  32'b00000001010001000000101111000011 ;
ROM[106] <=  32'b00001101010100010000101100001011 ;
ROM[107] <=  32'b00100100110101000100001100011101 ;
ROM[108] <=  32'b11010111011001010001000010010100 ;
ROM[109] <=  32'b01101100111000010100010000001110 ;
ROM[110] <=  32'b00110101001010110101000011110001 ;
ROM[111] <=  32'b11010110011001000001010000101100 ;
ROM[112] <=  32'b00000100000101101011010100001010 ;
ROM[113] <=  32'b00111101011011111010100101000010 ;
ROM[114] <=  32'b00000001111001010000011000000000 ;
ROM[115] <=  32'b00000000000000000000000000000000 ;
ROM[116] <=  32'b00000000000000000000000000000000 ;
ROM[117] <=  32'b00000000000000000000000000000001 ;
ROM[118] <=  32'b01000010100101101101011111101010 ;
ROM[119] <=  32'b01010001000000100000100000100001 ;
ROM[120] <=  32'b10010100010000101110000100101011 ;
ROM[121] <=  32'b01000101000100001011001100100110 ;
ROM[122] <=  32'b01000001010001000000011111001011 ;
ROM[123] <=  32'b00101000010100001011000101101000 ;
ROM[124] <=  32'b10001010000000000000000000000000 ;
ROM[125] <=  32'b00000000000001010000100100001001 ;
ROM[126] <=  32'b11010000010100010100000001100111 ;
ROM[127] <=  32'b10000010110111110000000000000000 ;
ROM[128] <=  32'b00000000000000000000000000000000 ;
ROM[129] <=  32'b00000000000000000000000000000000 ;
ROM[130] <=  32'b00000000000000000000000000000000 ;
ROM[131] <=  32'b00000000000000000000000000000000 ;
ROM[132] <=  32'b00000000000000000000000000000000 ;
ROM[133] <=  32'b00000000000000000000000000000000 ;
ROM[134] <=  32'b00000000000000000000000000000000 ;
ROM[135] <=  32'b00000000000000000000000000000000 ;
ROM[136] <=  32'b00000000000000000000000000000000 ;
ROM[137] <=  32'b00010100000100110110110001111110 ;
ROM[138] <=  32'b00110101000001010100100001101010 ;
ROM[139] <=  32'b10001100000000000000000000000000 ;
ROM[140] <=  32'b00000000000000000000000000000000 ;
ROM[141] <=  32'b00000000000000000000000000000000 ;
ROM[142] <=  32'b00000000000000000000000000000000 ;
ROM[143] <=  32'b00000000000000000000000000000000 ;
ROM[144] <=  32'b00000000000000000000000000000000 ;
ROM[145] <=  32'b00000000000000000000000000000000 ;
ROM[146] <=  32'b00000000000000000000000000000000 ;
ROM[147] <=  32'b00000000000000000000000101000000 ;
ROM[148] <=  32'b00010010010100100000011001010000 ;
ROM[149] <=  32'b01001000111111101110011010010100 ;
ROM[150] <=  32'b00011001101010000101101011110000 ;
ROM[151] <=  32'b00000000000000000000000000000000 ;
ROM[152] <=  32'b00000000000000000000000000000000 ;
ROM[153] <=  32'b00000000000000000000000000000000 ;
ROM[154] <=  32'b00000000000000000000000000000000 ;
ROM[155] <=  32'b00000101000001101001000011101000 ;
ROM[156] <=  32'b01110001010000110011011100001110 ;
ROM[157] <=  32'b10110100010100001110100001110111 ;
ROM[158] <=  32'b00000010000101000011101101001110 ;
ROM[159] <=  32'b10011100100001010000111010111110 ;
ROM[160] <=  32'b10011111111000010100001110000010 ;
ROM[161] <=  32'b11011100010011110101000010011111 ;
ROM[162] <=  32'b10001000001111101001001111001101 ;
ROM[163] <=  32'b00100000011101011111000000000000 ;
ROM[164] <=  32'b00000000000000000000000000000000 ;
ROM[165] <=  32'b00000000000000000000000000000000 ;
ROM[166] <=  32'b00000000000000000000000000010100 ;
ROM[167] <=  32'b00010010111110101111101000100101 ;
ROM[168] <=  32'b00001011101010110100010110111101 ;
ROM[169] <=  32'b01000011100010011000001101000001 ;
ROM[170] <=  32'b01010000110111011000010001111100 ;
ROM[171] <=  32'b10010100001100010111101000010110 ;
ROM[172] <=  32'b01100101000011100101011000000011 ;
ROM[173] <=  32'b10000001010000111011100000010011 ;
ROM[174] <=  32'b11010100010100001110110111101100 ;
ROM[175] <=  32'b01001111110101000011000101100100 ;
ROM[176] <=  32'b11001010010001001111111010111011 ;
ROM[177] <=  32'b11100010011100000000000000000000 ;
ROM[178] <=  32'b00000000000000000000000000000000 ;
ROM[179] <=  32'b00000000000000000001010000100111 ;
ROM[180] <=  32'b11110011110000000101010100000110 ;
ROM[181] <=  32'b11110100111000011001110000000000 ;
ROM[182] <=  32'b00000000000000000000000000000000 ;
ROM[183] <=  32'b00000000000000000000000000000000 ;
ROM[184] <=  32'b00000000000000000000000000000000 ;
ROM[185] <=  32'b00000000000000000000000000000000 ;
ROM[186] <=  32'b00000000000000000000000000000000 ;
ROM[187] <=  32'b01010000111010010111110001110010 ;
ROM[188] <=  32'b00010100001110010010110100101010 ;
ROM[189] <=  32'b10000101000010110100011110111111 ;
ROM[190] <=  32'b01100000000000000000000000000000 ;
ROM[191] <=  32'b00000000010100000100000010010101 ;
ROM[192] <=  32'b11101001110000000000000000000000 ;
ROM[193] <=  32'b00000000000000000000000000000000 ;
ROM[194] <=  32'b00000000000000000000000000000000 ;
ROM[195] <=  32'b00000000000000000000000000000000 ;
ROM[196] <=  32'b00000000000000000001010000101111 ;
ROM[197] <=  32'b01011000100100001110010100001100 ;
ROM[198] <=  32'b00011011000100100111000000000000 ;
ROM[199] <=  32'b00000000000000000000000000000000 ;
ROM[200] <=  32'b00000000000000000000000000010100 ;
ROM[201] <=  32'b00110100010101100101110111110101 ;
ROM[202] <=  32'b00001100111101010110010001110001 ;
ROM[203] <=  32'b01000000110011001100000101001111 ;
ROM[204] <=  32'b01010000010000100111101110010110 ;
ROM[205] <=  32'b10000000000000000000000000000000 ;
ROM[206] <=  32'b00000101000010100110011101000111 ;
ROM[207] <=  32'b10011101010000110101000000101011 ;
ROM[208] <=  32'b11101110010100001100111110000011 ;
ROM[209] <=  32'b10001111010101000010101101011001 ;
ROM[210] <=  32'b00011001010001010000110101000010 ;
ROM[211] <=  32'b01011101011111010100001011101110 ;
ROM[212] <=  32'b10101110001010000000000000000000 ;
ROM[213] <=  32'b00000000000000000001010000100000 ;
ROM[214] <=  32'b10100101110110000001010100001011 ;
ROM[215] <=  32'b10011100000010010000100101000010 ;
ROM[216] <=  32'b00100111101111111010111101010000 ;
ROM[217] <=  32'b01011110101011000000100010010100 ;
ROM[218] <=  32'b00101011010000111001111010110101 ;
ROM[219] <=  32'b00001010110000110100011011111001 ;
ROM[220] <=  32'b01000010101011111101011110101000 ;
ROM[221] <=  32'b01010000100010110101001110000100 ;
ROM[222] <=  32'b01000000000000000000000000000000 ;
ROM[223] <=  32'b00000101000010100010100101101000 ;
ROM[224] <=  32'b10100001010000110011000110010110 ;
ROM[225] <=  32'b11101000000000000000000000000000 ;
ROM[226] <=  32'b00000000000000000000000000000000 ;
ROM[227] <=  32'b00000000000001010000101101100111 ;
ROM[228] <=  32'b01110010110000010100001001000001 ;
ROM[229] <=  32'b00001010000000000000000000000000 ;
ROM[230] <=  32'b00000000000000000000000000000000 ;
ROM[231] <=  32'b00000000000000000000010100000110 ;
ROM[232] <=  32'b10101100110010110010110101000010 ;
ROM[233] <=  32'b11010110100110111100000101010000 ;
ROM[234] <=  32'b10110100111111000010100110000000 ;
ROM[235] <=  32'b00000000000000000000000000000000 ;
ROM[236] <=  32'b00000000000000000000000000000001 ;
ROM[237] <=  32'b01000010110000111000111101001011 ;
ROM[238] <=  32'b01010000101110111000011101000011 ;
ROM[239] <=  32'b00000000000000000000000000000000 ;
ROM[240] <=  32'b00000101000010010101010010010000 ;
ROM[241] <=  32'b00001001010000100101000111011010 ;
ROM[242] <=  32'b00110101010100001010100101010100 ;
ROM[243] <=  32'b01101101100000000000000000000000 ;
ROM[244] <=  32'b00000000000000000000000000000000 ;
ROM[245] <=  32'b00000000000000010100001101011110 ;
ROM[246] <=  32'b10000101011010000101000011100110 ;
ROM[247] <=  32'b01010000110011011001010000110000 ;
ROM[248] <=  32'b01111011000011010011010100001010 ;
ROM[249] <=  32'b01111111101101001011100101000011 ;
ROM[250] <=  32'b00001010101001110110111101010000 ;
ROM[251] <=  32'b11001101111011010101010000010100 ;
ROM[252] <=  32'b00100010101111100101011110110000 ;
ROM[253] <=  32'b00000000000000000000000000000001 ;
ROM[254] <=  32'b01000001100110010001111000001000 ;
ROM[255] <=  32'b01010000101001010100100000001000 ;
ROM[256] <=  32'b00010100001100000000111110000110 ;
ROM[257] <=  32'b01000000000000000000000000000000 ;
ROM[258] <=  32'b00000000000000000000000000000000 ;
ROM[259] <=  32'b00000000010100001110111000001001 ;
ROM[260] <=  32'b01111010000101000011110001011010 ;
ROM[261] <=  32'b10000100001101010000111010010101 ;
ROM[262] <=  32'b11011111011001010100001101100011 ;
ROM[263] <=  32'b11101101110100100101000010010000 ;
ROM[264] <=  32'b10100110011001111001010000100111 ;
ROM[265] <=  32'b10010111111110010001010011111110 ;
ROM[266] <=  32'b10100011110000100111000000000000 ;
ROM[267] <=  32'b00000000000000000000000001010000 ;
ROM[268] <=  32'b01000000010100100001101101010100 ;
ROM[269] <=  32'b00110001100010101010110001010101 ;
ROM[270] <=  32'b00001100001100110101101011011000 ;
ROM[271] <=  32'b00000000000000000000000000000000 ;
ROM[272] <=  32'b00000000000000000000000000000000 ;
ROM[273] <=  32'b00000000000000000000000000000000 ;
ROM[274] <=  32'b00000000000000000000000000000000 ;
ROM[275] <=  32'b00000000000000000000000000000000 ;
ROM[276] <=  32'b00000000000000000000000000000000 ;
ROM[277] <=  32'b00000000000000000000000000000000 ;
ROM[278] <=  32'b00000000000000000000000000000000 ;
ROM[279] <=  32'b00000000000000000000000000000000 ;
ROM[280] <=  32'b00000000000000000000000000000000 ;
ROM[281] <=  32'b00000000000000000001010000100011 ;
ROM[282] <=  32'b10011101111100011010010100001100 ;
ROM[283] <=  32'b10100000101011010011110101000011 ;
ROM[284] <=  32'b00010011001001000000111000000000 ;
ROM[285] <=  32'b00000000000000000000000000000000 ;
ROM[286] <=  32'b00000000000000000000000000000000 ;
ROM[287] <=  32'b00000000000000000000000000000001 ;
ROM[288] <=  32'b01000001110001010010111001100001 ;
ROM[289] <=  32'b01010000100011111001000111001101 ;
ROM[290] <=  32'b10010100000110101111100100101011 ;
ROM[291] <=  32'b10100000000000000000000000000000 ;
ROM[292] <=  32'b00000000000000000000000000000000 ;
ROM[293] <=  32'b00000000000000000000000000000000 ;
ROM[294] <=  32'b00000000000000000000000000000000 ;
ROM[295] <=  32'b00000000000001010000101100111111 ;
ROM[296] <=  32'b01110100101000010100001110000111 ;
ROM[297] <=  32'b00000011111110000101000011100101 ;
ROM[298] <=  32'b01010100101001100001010000111001 ;
ROM[299] <=  32'b11101101100010000001010100001101 ;
ROM[300] <=  32'b01110010111000010100100101000011 ;
ROM[301] <=  32'b00111110101100010000001001010000 ;
ROM[302] <=  32'b10011010001110100110001101000000 ;
ROM[303] <=  32'b00000000000000000000000000000000 ;
ROM[304] <=  32'b00000000000000000000000000000000 ;
ROM[305] <=  32'b00000000000000000000000000000000 ;
ROM[306] <=  32'b01001110110011101100010111001110 ;
ROM[307] <=  32'b01010011101100111011000101110011 ;
ROM[308] <=  32'b10010101000010000010011111001100 ;
ROM[309] <=  32'b00011001010000110011110110010001 ;
ROM[310] <=  32'b11010101010100001110011101100011 ;
ROM[311] <=  32'b01011110010101000011101100011011 ;
ROM[312] <=  32'b00010000101101010000111010011110 ;
ROM[313] <=  32'b00101111100011010100001100010001 ;
ROM[314] <=  32'b01001111100001000101000000001110 ;
ROM[315] <=  32'b00100100010101100101001110110011 ;
ROM[316] <=  32'b10110001011100111001010011101100 ;
ROM[317] <=  32'b11101100010111001110010100111011 ;
ROM[318] <=  32'b00111011000101110011100101001110 ;
ROM[319] <=  32'b11001110110001011100111001010100 ;
ROM[320] <=  32'b00011111001111110001101111110101 ;
ROM[321] <=  32'b00001110110001010110010001101101 ;
ROM[322] <=  32'b01000100000011111111010100010110 ;
ROM[323] <=  32'b01010001000100011101111110110111 ;
ROM[324] <=  32'b11010100010001111001111100000000 ;
ROM[325] <=  32'b10110101000100100010111011010010 ;
ROM[326] <=  32'b00100101010001001000001110001001 ;
ROM[327] <=  32'b11101011010100010000001111100110 ;
ROM[328] <=  32'b10110011110101000010101001111111 ;
ROM[329] <=  32'b00100101010101001110110011101100 ;
ROM[330] <=  32'b01011100111001010011101100111011 ;
ROM[331] <=  32'b00010111001110010100111011001110 ;
ROM[332] <=  32'b11000101110011100101010000110110 ;
ROM[333] <=  32'b11101011101110001100010100001111 ;
ROM[334] <=  32'b01010001010101101001000101000100 ;
ROM[335] <=  32'b00110101001111001001110101010001 ;
ROM[336] <=  32'b00100001101010101110100011010100 ;
ROM[337] <=  32'b01001001000000100001010101010101 ;
ROM[338] <=  32'b00010010101001110001101010010001 ;
ROM[339] <=  32'b01000100101101110001100001000000 ;
ROM[340] <=  32'b01010001001011011001110000011111 ;
ROM[341] <=  32'b10010100010000111101000001000001 ;
ROM[342] <=  32'b10010101000010111011011111011011 ;
ROM[343] <=  32'b10100001001110110011101100010111 ;
ROM[344] <=  32'b00111001010100000110001000010101 ;
ROM[345] <=  32'b01001000100101000011100111000101 ;
ROM[346] <=  32'b01101010100101010000111101001110 ;
ROM[347] <=  32'b10000011000110010100010001001011 ;
ROM[348] <=  32'b11000000110010110101000100011101 ;
ROM[349] <=  32'b10001001000101000101010001000101 ;
ROM[350] <=  32'b00010100110010001011010100010000 ;
ROM[351] <=  32'b11000010101110100000110101000100 ;
ROM[352] <=  32'b10010111010100111010000101010001 ;
ROM[353] <=  32'b00101101001101100010111110010100 ;
ROM[354] <=  32'b01001010111000100110000110010101 ;
ROM[355] <=  32'b00010000010010010010010001001101 ;
ROM[356] <=  32'b00111011001110110001011100111001 ;
ROM[357] <=  32'b01010000100110001111010101100000 ;
ROM[358] <=  32'b10010100001101110011001100010011 ;
ROM[359] <=  32'b01010101000100001001100101000110 ;
ROM[360] <=  32'b11111001010001000110010110001111 ;
ROM[361] <=  32'b00110100010100010000011101000100 ;
ROM[362] <=  32'b01001100100101000011111011010011 ;
ROM[363] <=  32'b11011000111001010000110000111011 ;
ROM[364] <=  32'b01111111110000010100001110100111 ;
ROM[365] <=  32'b10110010100101110101000100100100 ;
ROM[366] <=  32'b11111111100110110101010001001010 ;
ROM[367] <=  32'b11100100100111011111010100010001 ;
ROM[368] <=  32'b11000100011100110110110101000010 ;
ROM[369] <=  32'b11111010110000000000101001010000 ;
ROM[370] <=  32'b11000100010011000001001000010100 ;
ROM[371] <=  32'b00111000011100100001010111100101 ;
ROM[372] <=  32'b00010001110011101001010001110101 ;
ROM[373] <=  32'b01000100100011010111011110111011 ;
ROM[374] <=  32'b01010000111110001101101010001101 ;
ROM[375] <=  32'b01010100000110110011111110000101 ;
ROM[376] <=  32'b01010100111011001110110001011100 ;
ROM[377] <=  32'b11100100000000000000000000000000 ;
ROM[378] <=  32'b00000000010100010000010111100111 ;
ROM[379] <=  32'b00100000000101000100101000001010 ;
ROM[380] <=  32'b11100100000101010001001000101110 ;
ROM[381] <=  32'b00011011011001010100001110010000 ;
ROM[382] <=  32'b01100010001110100101000011000100 ;
ROM[383] <=  32'b11111000000100111101010000111011 ;
ROM[384] <=  32'b00110010011100001111010100010010 ;
ROM[385] <=  32'b01110000110000101101110101000100 ;
ROM[386] <=  32'b10010111100100000111010101010000 ;
ROM[387] <=  32'b11110110000011100000000111010011 ;
ROM[388] <=  32'b10110011101100010111001110010100 ;
ROM[389] <=  32'b11101100111011000101110011100101 ;
ROM[390] <=  32'b01000001110100111110110101000011 ;
ROM[391] <=  32'b01010000111000000011010001001110 ;
ROM[392] <=  32'b01010100010010001011010010110111 ;
ROM[393] <=  32'b11100101000100100011101110111000 ;
ROM[394] <=  32'b11100101010000111101001110110000 ;
ROM[395] <=  32'b00110111000000000000000000000000 ;
ROM[396] <=  32'b00000000000101000011100110100100 ;
ROM[397] <=  32'b01011001011001010001001010010100 ;
ROM[398] <=  32'b10010111001001010100010010111010 ;
ROM[399] <=  32'b00111000101100000101000100010001 ;
ROM[400] <=  32'b10010001011100001001010000101010 ;
ROM[401] <=  32'b10110110011100000011010100001010 ;
ROM[402] <=  32'b11111010110011101101000101000011 ;
ROM[403] <=  32'b10101111111101011011101101010000 ;
ROM[404] <=  32'b11101001000000001000100101010100 ;
ROM[405] <=  32'b01000100110100110100111101100101 ;
ROM[406] <=  32'b00010010001001011010001010101001 ;
ROM[407] <=  32'b01000011110100111011000010100001 ;
ROM[408] <=  32'b01001110110011101100010111001110 ;
ROM[409] <=  32'b01000000000000000000000000000000 ;
ROM[410] <=  32'b00000101000100011110000101011101 ;
ROM[411] <=  32'b11110101010001001011101000010101 ;
ROM[412] <=  32'b00010011010100010010110111011011 ;
ROM[413] <=  32'b10000101100101000100011100000101 ;
ROM[414] <=  32'b01110011100001010001000001111100 ;
ROM[415] <=  32'b00101100100110010100010000010011 ;
ROM[416] <=  32'b00101100001101100101000100001000 ;
ROM[417] <=  32'b01001111101110110101010001000111 ;
ROM[418] <=  32'b10100010101101101001010100010001 ;
ROM[419] <=  32'b10100000101110100000000101000011 ;
ROM[420] <=  32'b01001111101001011010111101001110 ;
ROM[421] <=  32'b11001110110001011100111001000000 ;
ROM[422] <=  32'b00000000000000000000000000000101 ;
ROM[423] <=  32'b00001101110001001001010001000101 ;
ROM[424] <=  32'b01000100100101000110100111101100 ;
ROM[425] <=  32'b01010001001011101010100100011101 ;
ROM[426] <=  32'b10010100010010101101100000010100 ;
ROM[427] <=  32'b11000101000100100100101011111011 ;
ROM[428] <=  32'b10001001010001000110011100100101 ;
ROM[429] <=  32'b10010010010100010001011111001110 ;
ROM[430] <=  32'b11011001000101000100011011101011 ;
ROM[431] <=  32'b11101001101001010001000010100100 ;
ROM[432] <=  32'b00010001001110010100000100100110 ;
ROM[433] <=  32'b10010000011000100100111011001110 ;
ROM[434] <=  32'b11000101110011100101001110110011 ;
ROM[435] <=  32'b10110001011100111001000000000000 ;
ROM[436] <=  32'b00000000000000000000000101000011 ;
ROM[437] <=  32'b01111001000101001001111101010001 ;
ROM[438] <=  32'b00011100001010110010110010010100 ;
ROM[439] <=  32'b01001000101000111010001101000101 ;
ROM[440] <=  32'b00010010001000011000010110000101 ;
ROM[441] <=  32'b01000100011000001110101010001010 ;
ROM[442] <=  32'b01010001000100100000110011001100 ;
ROM[443] <=  32'b01010100010000101111111110010011 ;
ROM[444] <=  32'b11100101000011010001000110010000 ;
ROM[445] <=  32'b11100001001110110011101100010111 ;
ROM[446] <=  32'b00111001010011101100111011000101 ;
ROM[447] <=  32'b11001110010100111011001110110001 ;
ROM[448] <=  32'b01110011100101001110110011101100 ;
ROM[449] <=  32'b01011100111001000000000000000000 ;
ROM[450] <=  32'b00000000000000000101000010001001 ;
ROM[451] <=  32'b10110101010001111001010000111001 ;
ROM[452] <=  32'b01101001101011101011010100001111 ;
ROM[453] <=  32'b10101111101111111010000101000011 ;
ROM[454] <=  32'b11101010100010100100000101010000 ;
ROM[455] <=  32'b11101001010001000000011110010100 ;
ROM[456] <=  32'b00110000001000111011110010000100 ;
ROM[457] <=  32'b11101100111011000101110011100101 ;
ROM[458] <=  32'b00111011001110110001011100111001 ;
ROM[459] <=  32'b01001110010110010001001111100110 ;
ROM[460] <=  32'b01010011100101100100010011111001 ;
ROM[461] <=  32'b10010101000010011011001001100000 ;
ROM[462] <=  32'b10101001010000111001101001011001 ;
ROM[463] <=  32'b00111000010100001111101000010011 ;
ROM[464] <=  32'b00001111000101000011111110010001 ;
ROM[465] <=  32'b11000001011001010000111011001111 ;
ROM[466] <=  32'b11011011000111010100001010100001 ;
ROM[467] <=  32'b10110000111110000000000000000000 ;
ROM[468] <=  32'b00000000000000000001001110010110 ;
ROM[469] <=  32'b01000100111110011001010011100101 ;
ROM[470] <=  32'b10010001001111100110010100111001 ;
ROM[471] <=  32'b01100100010011111001100101001110 ;
ROM[472] <=  32'b01011001000100111110011001010100 ;
ROM[473] <=  32'b00100101010001001100000111110101 ;
ROM[474] <=  32'b00010000000000001010001111001101 ;
ROM[475] <=  32'b01000100010000011101000001010001 ;
ROM[476] <=  32'b01010001000011110001000110001101 ;
ROM[477] <=  32'b11010100010000110001100000010100 ;
ROM[478] <=  32'b01110101000100000111011101011110 ;
ROM[479] <=  32'b10101001010000111101111000101000 ;
ROM[480] <=  32'b01110000010100001011100010111101 ;
ROM[481] <=  32'b00111111000000000000000000000000 ;
ROM[482] <=  32'b00000000000001001110010110010001 ;
ROM[483] <=  32'b00111110011001010011100101100100 ;
ROM[484] <=  32'b01001111100110010100111001011001 ;
ROM[485] <=  32'b00010011111001100101010000111100 ;
ROM[486] <=  32'b00000000111010010010010100010001 ;
ROM[487] <=  32'b10001110101101100000100101000100 ;
ROM[488] <=  32'b01110101001101100110010001010001 ;
ROM[489] <=  32'b00010101000101111111100001010100 ;
ROM[490] <=  32'b01000010100000100010001100100101 ;
ROM[491] <=  32'b00010000111111010000101010101001 ;
ROM[492] <=  32'b01000100010100011000110000001111 ;
ROM[493] <=  32'b01010001000001100101110000010011 ;
ROM[494] <=  32'b01000000000000000000000000000000 ;
ROM[495] <=  32'b00000000000000000000000000000000 ;
ROM[496] <=  32'b00000001001110010110010001001111 ;
ROM[497] <=  32'b10011001010100000111101101111010 ;
ROM[498] <=  32'b10111101000101000100001100101111 ;
ROM[499] <=  32'b01001011111101010001000111010001 ;
ROM[500] <=  32'b00101111000000010100010001001001 ;
ROM[501] <=  32'b00111001001011010101000100000000 ;
ROM[502] <=  32'b01100111111001111001010000111010 ;
ROM[503] <=  32'b01110000000001100111010100010000 ;
ROM[504] <=  32'b10101001010001001011100101000100 ;
ROM[505] <=  32'b01110110100100101001010001010001 ;
ROM[506] <=  32'b00011111101011011100110110010100 ;
ROM[507] <=  32'b00111101010110100100011000000000 ;
ROM[508] <=  32'b00000000000000000000000000000001 ;
ROM[509] <=  32'b00111001011001000100111110011001 ;
ROM[510] <=  32'b01010000101100001001010011100100 ;
ROM[511] <=  32'b01010100010001100000000110001111 ;
ROM[512] <=  32'b11000101000100100000101111111100 ;
ROM[513] <=  32'b10110101010000111011010111100100 ;
ROM[514] <=  32'b10101000010100001100010101110000 ;
ROM[515] <=  32'b11011101100101000011000101110000 ;
ROM[516] <=  32'b00101110110001010000111001010001 ;
ROM[517] <=  32'b10010100110010010100010001011101 ;
ROM[518] <=  32'b11001010111100000101000100100010 ;
ROM[519] <=  32'b00001010001100100101010001000100 ;
ROM[520] <=  32'b10111101100111111011000000000000 ;
ROM[521] <=  32'b00000000000000000000000100111001 ;
ROM[522] <=  32'b01100100010011111001100101010000 ;
ROM[523] <=  32'b11101101100101101111101010010100 ;
ROM[524] <=  32'b01000111110111110001010011010101 ;
ROM[525] <=  32'b00010010001010111001010001111001 ;
ROM[526] <=  32'b01000010110111101101100000010000 ;
ROM[527] <=  32'b01001111111110101100010000111100 ;
ROM[528] <=  32'b11010100000001111011111011010110 ;
ROM[529] <=  32'b10010101000010001001010001101000 ;
ROM[530] <=  32'b00111101010000111110101010001011 ;
ROM[531] <=  32'b10011110010100010010001011001011 ;
ROM[532] <=  32'b11101011100101000100100001110011 ;
ROM[533] <=  32'b11000000000001010000100010100001 ;
ROM[534] <=  32'b10100101110110000000000000000000 ;
ROM[535] <=  32'b00000000000000000101000011101110 ;
ROM[536] <=  32'b11111100111001101101010001001000 ;
ROM[537] <=  32'b00000100001001100111010100010010 ;
ROM[538] <=  32'b00100011010100100110100101000011 ;
ROM[539] <=  32'b00110100001101110001000100000000 ;
ROM[540] <=  32'b00000000000000000000000000010011 ;
ROM[541] <=  32'b10010110010001001111100110010100 ;
ROM[542] <=  32'b11100101100100010011111001100101 ;
ROM[543] <=  32'b01000011100001010010100001011011 ;
ROM[544] <=  32'b01010001000111100111010101011001 ;
ROM[545] <=  32'b10010100010010001101011000111100 ;
ROM[546] <=  32'b11100101000010100010010010111101 ;
ROM[547] <=  32'b01001100000000000000000000000000 ;
ROM[548] <=  32'b00000000010100001110011001110110 ;
ROM[549] <=  32'b11011010000101000100011111001011 ;
ROM[550] <=  32'b01011000100001010001001000111111 ;
ROM[551] <=  32'b01101101100011010100010000011101 ;
ROM[552] <=  32'b10100001110011110101000001010011 ;
ROM[553] <=  32'b00011101110101011101010000011000 ;
ROM[554] <=  32'b01000101100001100100010100001100 ;
ROM[555] <=  32'b10101010010110011111000101000100 ;
ROM[556] <=  32'b00011010011110101011111001010001 ;
ROM[557] <=  32'b00011111001001001111001000010100 ;
ROM[558] <=  32'b01000110101100001110100111000101 ;
ROM[559] <=  32'b00000101100000110111000011001100 ;
ROM[560] <=  32'b00000000000000000000000000000000 ;
ROM[561] <=  32'b01010000101100101110110001110001 ;
ROM[562] <=  32'b01010100010000011010000100110011 ;
ROM[563] <=  32'b11000101000100011110110101100001 ;
ROM[564] <=  32'b00100001010001000111001100101110 ;
ROM[565] <=  32'b10110101010100010000010000101010 ;
ROM[566] <=  32'b00000001010101000011110110110110 ;
ROM[567] <=  32'b11110110000001010001000000111101 ;
ROM[568] <=  32'b11110100100100010100010001010001 ;
ROM[569] <=  32'b10111010001001110101000100011011 ;
ROM[570] <=  32'b10001001010111111001010000111110 ;
ROM[571] <=  32'b00111111101001001011000000000000 ;
ROM[572] <=  32'b00000000000000000000000100111111 ;
ROM[573] <=  32'b10111000001011001101110101010000 ;
ROM[574] <=  32'b00100110101100101000000001010100 ;
ROM[575] <=  32'b00110110101000011110110111100101 ;
ROM[576] <=  32'b00010001010001100100000010011001 ;
ROM[577] <=  32'b01000100100000100110010101101110 ;
ROM[578] <=  32'b01010001000110011001011110101100 ;
ROM[579] <=  32'b11010100010001001000001111110101 ;
ROM[580] <=  32'b00100101000100001011001111110101 ;
ROM[581] <=  32'b10110001010001000011110111000101 ;
ROM[582] <=  32'b11001111010100010000010010000001 ;
ROM[583] <=  32'b00010100010101000001111110100101 ;
ROM[584] <=  32'b11001001110100000000000000000000 ;
ROM[585] <=  32'b00000000000000010011111111101001 ;
ROM[586] <=  32'b00100100010011100100111001011001 ;
ROM[587] <=  32'b00010011111001100101010000011101 ;
ROM[588] <=  32'b11011101101100101010010100001110 ;
ROM[589] <=  32'b01101011101101011101100101000100 ;
ROM[590] <=  32'b00101011100011110110100101010001 ;
ROM[591] <=  32'b00001111000101111001010111010100 ;
ROM[592] <=  32'b01000010101101110100100111010101 ;
ROM[593] <=  32'b00010000001011111011010000111001 ;
ROM[594] <=  32'b01000011110000001110100100000000 ;
ROM[595] <=  32'b01010000110011011111000110110000 ;
ROM[596] <=  32'b11010100000110110010001000011100 ;
ROM[597] <=  32'b11010101000001010011111011011000 ;
ROM[598] <=  32'b10111001001110010110010001001111 ;
ROM[599] <=  32'b10011001010011100101100100010011 ;
ROM[600] <=  32'b11100110010100111001011001000100 ;
ROM[601] <=  32'b11111001100101010000100111111100 ;
ROM[602] <=  32'b11010010110010010100001101010111 ;
ROM[603] <=  32'b00111010010111100101000011110000 ;
ROM[604] <=  32'b10111110101001100101010000111100 ;
ROM[605] <=  32'b11111000011100010010010100001110 ;
ROM[606] <=  32'b10000111110000011101010101000011 ;
ROM[607] <=  32'b01011101010000110010111001010000 ;
ROM[608] <=  32'b10101101010011001101010101010100 ;
ROM[609] <=  32'b00011100111100111111001111000100 ;
ROM[610] <=  32'b11100101100100010011111001100101 ;
ROM[611] <=  32'b00111001011001000100111110011001 ;
/*
ROM[1] <=  32'b00000000000000000000000000000000 ;
ROM[2] <=  32'b00000000000000000000000000000000 ;
ROM[3] <=  32'b00000101000010001001001010011000 ;
ROM[4] <=  32'b10010001010000110110101011101110 ;
ROM[5] <=  32'b10101011010100001110110101110001 ;
ROM[6] <=  32'b10100110010101000011110111111001 ;
ROM[7] <=  32'b10111001110001010000111110111111 ;
ROM[8] <=  32'b10111101111101010100001110010011 ;
ROM[9] <=  32'b00110010101001000101000010100001 ;
ROM[10] <=  32'b11010001111101010101010000000110 ;
ROM[11] <=  32'b00100011010010011010000000000000 ;
ROM[12] <=  32'b00000000000000000000000000000000 ;
ROM[13] <=  32'b00000000000000000000000000000000 ;
ROM[14] <=  32'b00000000000000000000000000010100 ;
ROM[15] <=  32'b00100000100101001010111111000101 ;
ROM[16] <=  32'b00001110010001100011001110101101 ;
ROM[17] <=  32'b01000100000000001110000111010010 ;
ROM[18] <=  32'b01010001000001011001001001011110 ;
ROM[19] <=  32'b11010100010000101000111100001111 ;
ROM[20] <=  32'b11100101000100001100010110010100 ;
ROM[21] <=  32'b10101101010001000011000011101011 ;
ROM[22] <=  32'b11000110010100010000010011001011 ;
ROM[23] <=  32'b10010111110101000011001011110101 ;
ROM[24] <=  32'b10000000000101010000010111110011 ;
ROM[25] <=  32'b00001000100011000000000000000000 ;
ROM[26] <=  32'b00000000000000000000000000000000 ;
ROM[27] <=  32'b00000000000000000001010000110100 ;
ROM[28] <=  32'b11001111111100000010010100001110 ;
ROM[29] <=  32'b01101000000000000110000101000011 ;
ROM[30] <=  32'b11010001010101101111111101010000 ;
ROM[31] <=  32'b11110101110000101000011001010100 ;
ROM[32] <=  32'b00110101000010011111111011010101 ;
ROM[33] <=  32'b00001110111110010011001111001001 ;
ROM[34] <=  32'b01000100000111100100011110100010 ;
ROM[35] <=  32'b01010001000010011101010010010000 ;
ROM[36] <=  32'b10010100001111111110001111010010 ;
ROM[37] <=  32'b10010101000011001010110010011101 ;
ROM[38] <=  32'b01010000000000000000000000000000 ;
ROM[39] <=  32'b00000000010100000110100000100000 ;
ROM[40] <=  32'b00010110010101000011010000100000 ;
ROM[41] <=  32'b11110100000001010000110110110011 ;
ROM[42] <=  32'b11100111100010010100001011011010 ;
ROM[43] <=  32'b01111101000001110000000000000000 ;
ROM[44] <=  32'b00000000000000000000000000000000 ;
ROM[45] <=  32'b00000000000000000000000000000000 ;
ROM[46] <=  32'b00000000000000000000000101000001 ;
ROM[47] <=  32'b01011111111101110101110101010000 ;
ROM[48] <=  32'b11111101011000011111011100010100 ;
ROM[49] <=  32'b00111111111011100100101010000101 ;
ROM[50] <=  32'b00001110100111000010100110011101 ;
ROM[51] <=  32'b01000010000101101110111111110100 ;
ROM[52] <=  32'b01010000100011010001110110010011 ;
ROM[53] <=  32'b10010100001100000100110100010010 ;
ROM[54] <=  32'b11110101000011001000001000110010 ;
ROM[55] <=  32'b10011101010000101011101101101010 ;
ROM[56] <=  32'b11110110010100000101000011110100 ;
ROM[57] <=  32'b10100101000000000000000000000000 ;
ROM[58] <=  32'b00000000000001010000001111001111 ;
ROM[59] <=  32'b11110101000000000000000000000000 ;
ROM[60] <=  32'b00000000000000000101000010110010 ;
ROM[61] <=  32'b10001111000011100001010000111011 ;
ROM[62] <=  32'b11011110111111000011010100001110 ;
ROM[63] <=  32'b11011000110000011110000101000010 ;
ROM[64] <=  32'b11011101111001101110111001010000 ;
ROM[65] <=  32'b10111111010010110011100101010100 ;
ROM[66] <=  32'b00110001111001110111001011100101 ;
ROM[67] <=  32'b00001100110011010001010000111101 ;
ROM[68] <=  32'b01000011011000110010001100011100 ;
ROM[69] <=  32'b01010000110011001101110011111111 ;
ROM[70] <=  32'b10010100000011111111000101000101 ;
ROM[71] <=  32'b01010000000000000000000000000000 ;
ROM[72] <=  32'b00000000000000000000000000000000 ;
ROM[73] <=  32'b00000000000000000000000000000000 ;
ROM[74] <=  32'b00000000000101000011100010100111 ;
ROM[75] <=  32'b10011011110001010000111001110010 ;
ROM[76] <=  32'b00001101000010010100001100111010 ;
ROM[77] <=  32'b10010111111000000101000010100010 ;
ROM[78] <=  32'b10101100001111111101010000110001 ;
ROM[79] <=  32'b01101010000100010101010100001110 ;
ROM[80] <=  32'b00110010111111000011100101000011 ;
ROM[81] <=  32'b10100001011101101001111101010000 ;
ROM[82] <=  32'b11010100010010000110011111010011 ;
ROM[83] <=  32'b11111001111100011100001000110000 ;
ROM[84] <=  32'b00000000000000000000000000000001 ;
ROM[85] <=  32'b01000010011001011000110111000110 ;
ROM[86] <=  32'b01010000100101100111110001101011 ;
ROM[87] <=  32'b00010100001100011100001110001110 ;
ROM[88] <=  32'b00110101000011100010010111011101 ;
ROM[89] <=  32'b01011001010000110011111000111001 ;
ROM[90] <=  32'b11001111000000000000000000000000 ;
ROM[91] <=  32'b00000000000000000000000000000000 ;
ROM[92] <=  32'b00000000000001010000111001001010 ;
ROM[93] <=  32'b11110011010010010100010000010000 ;
ROM[94] <=  32'b00111110000011100101000100000010 ;
ROM[95] <=  32'b00110011000000111001010000110010 ;
ROM[96] <=  32'b11010011101101001011010100001100 ;
ROM[97] <=  32'b00001101110011011001010101000011 ;
ROM[98] <=  32'b10010101111110100011001101010000 ;
ROM[99] <=  32'b11100010101110100011011001010100 ;
ROM[100] <=  32'b00101000111100011110001000100101 ;
ROM[101] <=  32'b00001100011010111010011100001101 ;
ROM[102] <=  32'b01000011000010001011110000110010 ;
ROM[103] <=  32'b00000000000000000000000000000000 ;
ROM[104] <=  32'b00000000000000000000000000000000 ;
ROM[105] <=  32'b00000000000000000000000000000000 ;
ROM[106] <=  32'b00000001010001000000101111000011 ;
ROM[107] <=  32'b00001101010100010000101100001011 ;
ROM[108] <=  32'b00100100110101000100001100011101 ;
ROM[109] <=  32'b11010111011001010001000010010100 ;
ROM[110] <=  32'b01101100111000010100010000001110 ;
ROM[111] <=  32'b00110101001010110101000011110001 ;
ROM[112] <=  32'b11010110011001000001010000101100 ;
ROM[113] <=  32'b00000100000101101011010100001010 ;
ROM[114] <=  32'b00111101011011111010100101000010 ;
ROM[115] <=  32'b00000001111001010000011000000000 ;
ROM[116] <=  32'b00000000000000000000000000000000 ;
ROM[117] <=  32'b00000000000000000000000000000000 ;
ROM[118] <=  32'b00000000000000000000000000000001 ;
ROM[119] <=  32'b01000010100101101101011111101010 ;
ROM[120] <=  32'b01010001000000100000100000100001 ;
ROM[121] <=  32'b10010100010000101110000100101011 ;
ROM[122] <=  32'b01000101000100001011001100100110 ;
ROM[123] <=  32'b01000001010001000000011111001011 ;
ROM[124] <=  32'b00101000010100001011000101101000 ;
ROM[125] <=  32'b10001010000000000000000000000000 ;
ROM[126] <=  32'b00000000000001010000100100001001 ;
ROM[127] <=  32'b11010000010100010100000001100111 ;
ROM[128] <=  32'b10000010110111110000000000000000 ;
ROM[129] <=  32'b00000000000000000000000000000000 ;
ROM[130] <=  32'b00000000000000000000000000000000 ;
ROM[131] <=  32'b00000000000000000000000000000000 ;
ROM[132] <=  32'b00000000000000000000000000000000 ;
ROM[133] <=  32'b00000000000000000000000000000000 ;
ROM[134] <=  32'b00000000000000000000000000000000 ;
ROM[135] <=  32'b00000000000000000000000000000000 ;
ROM[136] <=  32'b00000000000000000000000000000000 ;
ROM[137] <=  32'b00000000000000000000000000000000 ;
ROM[138] <=  32'b00010100000100110110110001111110 ;
ROM[139] <=  32'b00110101000001010100100001101010 ;
ROM[140] <=  32'b10001100000000000000000000000000 ;
ROM[141] <=  32'b00000000000000000000000000000000 ;
ROM[142] <=  32'b00000000000000000000000000000000 ;
ROM[143] <=  32'b00000000000000000000000000000000 ;
ROM[144] <=  32'b00000000000000000000000000000000 ;
ROM[145] <=  32'b00000000000000000000000000000000 ;
ROM[146] <=  32'b00000000000000000000000000000000 ;
ROM[147] <=  32'b00000000000000000000000000000000 ;
ROM[148] <=  32'b00000000000000000000000101000000 ;
ROM[149] <=  32'b00010010010100100000011001010000 ;
ROM[150] <=  32'b01001000111111101110011010010100 ;
ROM[151] <=  32'b00011001101010000101101011110000 ;
ROM[152] <=  32'b00000000000000000000000000000000 ;
ROM[153] <=  32'b00000000000000000000000000000000 ;
ROM[154] <=  32'b00000000000000000000000000000000 ;
ROM[155] <=  32'b00000000000000000000000000000000 ;
ROM[156] <=  32'b00000101000001101001000011101000 ;
ROM[157] <=  32'b01110001010000110011011100001110 ;
ROM[158] <=  32'b10110100010100001110100001110111 ;
ROM[159] <=  32'b00000010000101000011101101001110 ;
ROM[160] <=  32'b10011100100001010000111010111110 ;
ROM[161] <=  32'b10011111111000010100001110000010 ;
ROM[162] <=  32'b11011100010011110101000010011111 ;
ROM[163] <=  32'b10001000001111101001001111001101 ;
ROM[164] <=  32'b00100000011101011111000000000000 ;
ROM[165] <=  32'b00000000000000000000000000000000 ;
ROM[166] <=  32'b00000000000000000000000000000000 ;
ROM[167] <=  32'b00000000000000000000000000010100 ;
ROM[168] <=  32'b00010010111110101111101000100101 ;
ROM[169] <=  32'b00001011101010110100010110111101 ;
ROM[170] <=  32'b01000011100010011000001101000001 ;
ROM[171] <=  32'b01010000110111011000010001111100 ;
ROM[172] <=  32'b10010100001100010111101000010110 ;
ROM[173] <=  32'b01100101000011100101011000000011 ;
ROM[174] <=  32'b10000001010000111011100000010011 ;
ROM[175] <=  32'b11010100010100001110110111101100 ;
ROM[176] <=  32'b01001111110101000011000101100100 ;
ROM[177] <=  32'b11001010010001001111111010111011 ;
ROM[178] <=  32'b11100010011100000000000000000000 ;
ROM[179] <=  32'b00000000000000000000000000000000 ;
ROM[180] <=  32'b00000000000000000001010000100111 ;
ROM[181] <=  32'b11110011110000000101010100000110 ;
ROM[182] <=  32'b11110100111000011001110000000000 ;
ROM[183] <=  32'b00000000000000000000000000000000 ;
ROM[184] <=  32'b00000000000000000000000000000000 ;
ROM[185] <=  32'b00000000000000000000000000000000 ;
ROM[186] <=  32'b00000000000000000000000000000000 ;
ROM[187] <=  32'b00000000000000000000000000000000 ;
ROM[188] <=  32'b01010000111010010111110001110010 ;
ROM[189] <=  32'b00010100001110010010110100101010 ;
ROM[190] <=  32'b10000101000010110100011110111111 ;
ROM[191] <=  32'b01100000000000000000000000000000 ;
ROM[192] <=  32'b00000000010100000100000010010101 ;
ROM[193] <=  32'b11101001110000000000000000000000 ;
ROM[194] <=  32'b00000000000000000000000000000000 ;
ROM[195] <=  32'b00000000000000000000000000000000 ;
ROM[196] <=  32'b00000000000000000000000000000000 ;
ROM[197] <=  32'b00000000000000000001010000101111 ;
ROM[198] <=  32'b01011000100100001110010100001100 ;
ROM[199] <=  32'b00011011000100100111000000000000 ;
ROM[200] <=  32'b00000000000000000000000000000000 ;
ROM[201] <=  32'b00000000000000000000000000010100 ;
ROM[202] <=  32'b00110100010101100101110111110101 ;
ROM[203] <=  32'b00001100111101010110010001110001 ;
ROM[204] <=  32'b01000000110011001100000101001111 ;
ROM[205] <=  32'b01010000010000100111101110010110 ;
ROM[206] <=  32'b10000000000000000000000000000000 ;
ROM[207] <=  32'b00000101000010100110011101000111 ;
ROM[208] <=  32'b10011101010000110101000000101011 ;
ROM[209] <=  32'b11101110010100001100111110000011 ;
ROM[210] <=  32'b10001111010101000010101101011001 ;
ROM[211] <=  32'b00011001010001010000110101000010 ;
ROM[212] <=  32'b01011101011111010100001011101110 ;
ROM[213] <=  32'b10101110001010000000000000000000 ;
ROM[214] <=  32'b00000000000000000001010000100000 ;
ROM[215] <=  32'b10100101110110000001010100001011 ;
ROM[216] <=  32'b10011100000010010000100101000010 ;
ROM[217] <=  32'b00100111101111111010111101010000 ;
ROM[218] <=  32'b01011110101011000000100010010100 ;
ROM[219] <=  32'b00101011010000111001111010110101 ;
ROM[220] <=  32'b00001010110000110100011011111001 ;
ROM[221] <=  32'b01000010101011111101011110101000 ;
ROM[222] <=  32'b01010000100010110101001110000100 ;
ROM[223] <=  32'b01000000000000000000000000000000 ;
ROM[224] <=  32'b00000101000010100010100101101000 ;
ROM[225] <=  32'b10100001010000110011000110010110 ;
ROM[226] <=  32'b11101000000000000000000000000000 ;
ROM[227] <=  32'b00000000000000000000000000000000 ;
ROM[228] <=  32'b00000000000001010000101101100111 ;
ROM[229] <=  32'b01110010110000010100001001000001 ;
ROM[230] <=  32'b00001010000000000000000000000000 ;
ROM[231] <=  32'b00000000000000000000000000000000 ;
ROM[232] <=  32'b00000000000000000000010100000110 ;
ROM[233] <=  32'b10101100110010110010110101000010 ;
ROM[234] <=  32'b11010110100110111100000101010000 ;
ROM[235] <=  32'b10110100111111000010100110000000 ;
ROM[236] <=  32'b00000000000000000000000000000000 ;
ROM[237] <=  32'b00000000000000000000000000000001 ;
ROM[238] <=  32'b01000010110000111000111101001011 ;
ROM[239] <=  32'b01010000101110111000011101000011 ;
ROM[240] <=  32'b00000000000000000000000000000000 ;
ROM[241] <=  32'b00000101000010010101010010010000 ;
ROM[242] <=  32'b00001001010000100101000111011010 ;
ROM[243] <=  32'b00110101010100001010100101010100 ;
ROM[244] <=  32'b01101101100000000000000000000000 ;
ROM[245] <=  32'b00000000000000000000000000000000 ;
ROM[246] <=  32'b00000000000000010100001101011110 ;
ROM[247] <=  32'b10000101011010000101000011100110 ;
ROM[248] <=  32'b01010000110011011001010000110000 ;
ROM[249] <=  32'b01111011000011010011010100001010 ;
ROM[250] <=  32'b01111111101101001011100101000011 ;
ROM[251] <=  32'b00001010101001110110111101010000 ;
ROM[252] <=  32'b11001101111011010101010000010100 ;
ROM[253] <=  32'b00100010101111100101011110110000 ;
ROM[254] <=  32'b00000000000000000000000000000001 ;
ROM[255] <=  32'b01000001100110010001111000001000 ;
ROM[256] <=  32'b01010000101001010100100000001000 ;
ROM[257] <=  32'b00010100001100000000111110000110 ;
ROM[258] <=  32'b01000000000000000000000000000000 ;
ROM[259] <=  32'b00000000000000000000000000000000 ;
ROM[260] <=  32'b00000000010100001110111000001001 ;
ROM[261] <=  32'b01111010000101000011110001011010 ;
ROM[262] <=  32'b10000100001101010000111010010101 ;
ROM[263] <=  32'b11011111011001010100001101100011 ;
ROM[264] <=  32'b11101101110100100101000010010000 ;
ROM[265] <=  32'b10100110011001111001010000100111 ;
ROM[266] <=  32'b10010111111110010001010011111110 ;
ROM[267] <=  32'b10100011110000100111000000000000 ;
ROM[268] <=  32'b00000000000000000000000001010000 ;
ROM[269] <=  32'b01000000010100100001101101010100 ;
ROM[270] <=  32'b00110001100010101010110001010101 ;
ROM[271] <=  32'b00001100001100110101101011011000 ;
ROM[272] <=  32'b00000000000000000000000000000000 ;
ROM[273] <=  32'b00000000000000000000000000000000 ;
ROM[274] <=  32'b00000000000000000000000000000000 ;
ROM[275] <=  32'b00000000000000000000000000000000 ;
ROM[276] <=  32'b00000000000000000000000000000000 ;
ROM[277] <=  32'b00000000000000000000000000000000 ;
ROM[278] <=  32'b00000000000000000000000000000000 ;
ROM[279] <=  32'b00000000000000000000000000000000 ;
ROM[280] <=  32'b00000000000000000000000000000000 ;
ROM[281] <=  32'b00000000000000000000000000000000 ;
ROM[282] <=  32'b00000000000000000001010000100011 ;
ROM[283] <=  32'b10011101111100011010010100001100 ;
ROM[284] <=  32'b10100000101011010011110101000011 ;
ROM[285] <=  32'b00010011001001000000111000000000 ;
ROM[286] <=  32'b00000000000000000000000000000000 ;
ROM[287] <=  32'b00000000000000000000000000000000 ;
ROM[288] <=  32'b00000000000000000000000000000001 ;
ROM[289] <=  32'b01000001110001010010111001100001 ;
ROM[290] <=  32'b01010000100011111001000111001101 ;
ROM[291] <=  32'b10010100000110101111100100101011 ;
ROM[292] <=  32'b10100000000000000000000000000000 ;
ROM[293] <=  32'b00000000000000000000000000000000 ;
ROM[294] <=  32'b00000000000000000000000000000000 ;
ROM[295] <=  32'b00000000000000000000000000000000 ;
ROM[296] <=  32'b00000000000001010000101100111111 ;
ROM[297] <=  32'b01110100101000010100001110000111 ;
ROM[298] <=  32'b00000011111110000101000011100101 ;
ROM[299] <=  32'b01010100101001100001010000111001 ;
ROM[300] <=  32'b11101101100010000001010100001101 ;
ROM[301] <=  32'b01110010111000010100100101000011 ;
ROM[302] <=  32'b00111110101100010000001001010000 ;
ROM[303] <=  32'b10011010001110100110001101000000 ;
ROM[304] <=  32'b00000000000000000000000000000000 ;
ROM[305] <=  32'b00000000000000000000000000000000 ;
ROM[306] <=  32'b00000000000000000000000000000000 ;
ROM[307] <=  32'b01001110110011101100010111001110 ;
ROM[308] <=  32'b01010011101100111011000101110011 ;
ROM[309] <=  32'b10010101000010000010011111001100 ;
ROM[310] <=  32'b00011001010000110011110110010001 ;
ROM[311] <=  32'b11010101010100001110011101100011 ;
ROM[312] <=  32'b01011110010101000011101100011011 ;
ROM[313] <=  32'b00010000101101010000111010011110 ;
ROM[314] <=  32'b00101111100011010100001100010001 ;
ROM[315] <=  32'b01001111100001000101000000001110 ;
ROM[316] <=  32'b00100100010101100101001110110011 ;
ROM[317] <=  32'b10110001011100111001010011101100 ;
ROM[318] <=  32'b11101100010111001110010100111011 ;
ROM[319] <=  32'b00111011000101110011100101001110 ;
ROM[320] <=  32'b11001110110001011100111001010100 ;
ROM[321] <=  32'b00011111001111110001101111110101 ;
ROM[322] <=  32'b00001110110001010110010001101101 ;
ROM[323] <=  32'b01000100000011111111010100010110 ;
ROM[324] <=  32'b01010001000100011101111110110111 ;
ROM[325] <=  32'b11010100010001111001111100000000 ;
ROM[326] <=  32'b10110101000100100010111011010010 ;
ROM[327] <=  32'b00100101010001001000001110001001 ;
ROM[328] <=  32'b11101011010100010000001111100110 ;
ROM[329] <=  32'b10110011110101000010101001111111 ;
ROM[330] <=  32'b00100101010101001110110011101100 ;
ROM[331] <=  32'b01011100111001010011101100111011 ;
ROM[332] <=  32'b00010111001110010100111011001110 ;
ROM[333] <=  32'b11000101110011100101010000110110 ;
ROM[334] <=  32'b11101011101110001100010100001111 ;
ROM[335] <=  32'b01010001010101101001000101000100 ;
ROM[336] <=  32'b00110101001111001001110101010001 ;
ROM[337] <=  32'b00100001101010101110100011010100 ;
ROM[338] <=  32'b01001001000000100001010101010101 ;
ROM[339] <=  32'b00010010101001110001101010010001 ;
ROM[340] <=  32'b01000100101101110001100001000000 ;
ROM[341] <=  32'b01010001001011011001110000011111 ;
ROM[342] <=  32'b10010100010000111101000001000001 ;
ROM[343] <=  32'b10010101000010111011011111011011 ;
ROM[344] <=  32'b10100001001110110011101100010111 ;
ROM[345] <=  32'b00111001010100000110001000010101 ;
ROM[346] <=  32'b01001000100101000011100111000101 ;
ROM[347] <=  32'b01101010100101010000111101001110 ;
ROM[348] <=  32'b10000011000110010100010001001011 ;
ROM[349] <=  32'b11000000110010110101000100011101 ;
ROM[350] <=  32'b10001001000101000101010001000101 ;
ROM[351] <=  32'b00010100110010001011010100010000 ;
ROM[352] <=  32'b11000010101110100000110101000100 ;
ROM[353] <=  32'b10010111010100111010000101010001 ;
ROM[354] <=  32'b00101101001101100010111110010100 ;
ROM[355] <=  32'b01001010111000100110000110010101 ;
ROM[356] <=  32'b00010000010010010010010001001101 ;
ROM[357] <=  32'b00111011001110110001011100111001 ;
ROM[358] <=  32'b01010000100110001111010101100000 ;
ROM[359] <=  32'b10010100001101110011001100010011 ;
ROM[360] <=  32'b01010101000100001001100101000110 ;
ROM[361] <=  32'b11111001010001000110010110001111 ;
ROM[362] <=  32'b00110100010100010000011101000100 ;
ROM[363] <=  32'b01001100100101000011111011010011 ;
ROM[364] <=  32'b11011000111001010000110000111011 ;
ROM[365] <=  32'b01111111110000010100001110100111 ;
ROM[366] <=  32'b10110010100101110101000100100100 ;
ROM[367] <=  32'b11111111100110110101010001001010 ;
ROM[368] <=  32'b11100100100111011111010100010001 ;
ROM[369] <=  32'b11000100011100110110110101000010 ;
ROM[370] <=  32'b11111010110000000000101001010000 ;
ROM[371] <=  32'b11000100010011000001001000010100 ;
ROM[372] <=  32'b00111000011100100001010111100101 ;
ROM[373] <=  32'b00010001110011101001010001110101 ;
ROM[374] <=  32'b01000100100011010111011110111011 ;
ROM[375] <=  32'b01010000111110001101101010001101 ;
ROM[376] <=  32'b01010100000110110011111110000101 ;
ROM[377] <=  32'b01010100111011001110110001011100 ;
ROM[378] <=  32'b11100100000000000000000000000000 ;
ROM[379] <=  32'b00000000010100010000010111100111 ;
ROM[380] <=  32'b00100000000101000100101000001010 ;
ROM[381] <=  32'b11100100000101010001001000101110 ;
ROM[382] <=  32'b00011011011001010100001110010000 ;
ROM[383] <=  32'b01100010001110100101000011000100 ;
ROM[384] <=  32'b11111000000100111101010000111011 ;
ROM[385] <=  32'b00110010011100001111010100010010 ;
ROM[386] <=  32'b01110000110000101101110101000100 ;
ROM[387] <=  32'b10010111100100000111010101010000 ;
ROM[388] <=  32'b11110110000011100000000111010011 ;
ROM[389] <=  32'b10110011101100010111001110010100 ;
ROM[390] <=  32'b11101100111011000101110011100101 ;
ROM[391] <=  32'b01000001110100111110110101000011 ;
ROM[392] <=  32'b01010000111000000011010001001110 ;
ROM[393] <=  32'b01010100010010001011010010110111 ;
ROM[394] <=  32'b11100101000100100011101110111000 ;
ROM[395] <=  32'b11100101010000111101001110110000 ;
ROM[396] <=  32'b00110111000000000000000000000000 ;
ROM[397] <=  32'b00000000000101000011100110100100 ;
ROM[398] <=  32'b01011001011001010001001010010100 ;
ROM[399] <=  32'b10010111001001010100010010111010 ;
ROM[400] <=  32'b00111000101100000101000100010001 ;
ROM[401] <=  32'b10010001011100001001010000101010 ;
ROM[402] <=  32'b10110110011100000011010100001010 ;
ROM[403] <=  32'b11111010110011101101000101000011 ;
ROM[404] <=  32'b10101111111101011011101101010000 ;
ROM[405] <=  32'b11101001000000001000100101010100 ;
ROM[406] <=  32'b01000100110100110100111101100101 ;
ROM[407] <=  32'b00010010001001011010001010101001 ;
ROM[408] <=  32'b01000011110100111011000010100001 ;
ROM[409] <=  32'b01001110110011101100010111001110 ;
ROM[410] <=  32'b01000000000000000000000000000000 ;
ROM[411] <=  32'b00000101000100011110000101011101 ;
ROM[412] <=  32'b11110101010001001011101000010101 ;
ROM[413] <=  32'b00010011010100010010110111011011 ;
ROM[414] <=  32'b10000101100101000100011100000101 ;
ROM[415] <=  32'b01110011100001010001000001111100 ;
ROM[416] <=  32'b00101100100110010100010000010011 ;
ROM[417] <=  32'b00101100001101100101000100001000 ;
ROM[418] <=  32'b01001111101110110101010001000111 ;
ROM[419] <=  32'b10100010101101101001010100010001 ;
ROM[420] <=  32'b10100000101110100000000101000011 ;
ROM[421] <=  32'b01001111101001011010111101001110 ;
ROM[422] <=  32'b11001110110001011100111001000000 ;
ROM[423] <=  32'b00000000000000000000000000000101 ;
ROM[424] <=  32'b00001101110001001001010001000101 ;
ROM[425] <=  32'b01000100100101000110100111101100 ;
ROM[426] <=  32'b01010001001011101010100100011101 ;
ROM[427] <=  32'b10010100010010101101100000010100 ;
ROM[428] <=  32'b11000101000100100100101011111011 ;
ROM[429] <=  32'b10001001010001000110011100100101 ;
ROM[430] <=  32'b10010010010100010001011111001110 ;
ROM[431] <=  32'b11011001000101000100011011101011 ;
ROM[432] <=  32'b11101001101001010001000010100100 ;
ROM[433] <=  32'b00010001001110010100000100100110 ;
ROM[434] <=  32'b10010000011000100100111011001110 ;
ROM[435] <=  32'b11000101110011100101001110110011 ;
ROM[436] <=  32'b10110001011100111001000000000000 ;
ROM[437] <=  32'b00000000000000000000000101000011 ;
ROM[438] <=  32'b01111001000101001001111101010001 ;
ROM[439] <=  32'b00011100001010110010110010010100 ;
ROM[440] <=  32'b01001000101000111010001101000101 ;
ROM[441] <=  32'b00010010001000011000010110000101 ;
ROM[442] <=  32'b01000100011000001110101010001010 ;
ROM[443] <=  32'b01010001000100100000110011001100 ;
ROM[444] <=  32'b01010100010000101111111110010011 ;
ROM[445] <=  32'b11100101000011010001000110010000 ;
ROM[446] <=  32'b11100001001110110011101100010111 ;
ROM[447] <=  32'b00111001010011101100111011000101 ;
ROM[448] <=  32'b11001110010100111011001110110001 ;
ROM[449] <=  32'b01110011100101001110110011101100 ;
ROM[450] <=  32'b01011100111001000000000000000000 ;
ROM[451] <=  32'b00000000000000000101000010001001 ;
ROM[452] <=  32'b10110101010001111001010000111001 ;
ROM[453] <=  32'b01101001101011101011010100001111 ;
ROM[454] <=  32'b10101111101111111010000101000011 ;
ROM[455] <=  32'b11101010100010100100000101010000 ;
ROM[456] <=  32'b11101001010001000000011110010100 ;
ROM[457] <=  32'b00110000001000111011110010000100 ;
ROM[458] <=  32'b11101100111011000101110011100101 ;
ROM[459] <=  32'b00111011001110110001011100111001 ;
ROM[460] <=  32'b01001110010110010001001111100110 ;
ROM[461] <=  32'b01010011100101100100010011111001 ;
ROM[462] <=  32'b10010101000010011011001001100000 ;
ROM[463] <=  32'b10101001010000111001101001011001 ;
ROM[464] <=  32'b00111000010100001111101000010011 ;
ROM[465] <=  32'b00001111000101000011111110010001 ;
ROM[466] <=  32'b11000001011001010000111011001111 ;
ROM[467] <=  32'b11011011000111010100001010100001 ;
ROM[468] <=  32'b10110000111110000000000000000000 ;
ROM[469] <=  32'b00000000000000000001001110010110 ;
ROM[470] <=  32'b01000100111110011001010011100101 ;
ROM[471] <=  32'b10010001001111100110010100111001 ;
ROM[472] <=  32'b01100100010011111001100101001110 ;
ROM[473] <=  32'b01011001000100111110011001010100 ;
ROM[474] <=  32'b00100101010001001100000111110101 ;
ROM[475] <=  32'b00010000000000001010001111001101 ;
ROM[476] <=  32'b01000100010000011101000001010001 ;
ROM[477] <=  32'b01010001000011110001000110001101 ;
ROM[478] <=  32'b11010100010000110001100000010100 ;
ROM[479] <=  32'b01110101000100000111011101011110 ;
ROM[480] <=  32'b10101001010000111101111000101000 ;
ROM[481] <=  32'b01110000010100001011100010111101 ;
ROM[482] <=  32'b00111111000000000000000000000000 ;
ROM[483] <=  32'b00000000000001001110010110010001 ;
ROM[484] <=  32'b00111110011001010011100101100100 ;
ROM[485] <=  32'b01001111100110010100111001011001 ;
ROM[486] <=  32'b00010011111001100101010000111100 ;
ROM[487] <=  32'b00000000111010010010010100010001 ;
ROM[488] <=  32'b10001110101101100000100101000100 ;
ROM[489] <=  32'b01110101001101100110010001010001 ;
ROM[490] <=  32'b00010101000101111111100001010100 ;
ROM[491] <=  32'b01000010100000100010001100100101 ;
ROM[492] <=  32'b00010000111111010000101010101001 ;
ROM[493] <=  32'b01000100010100011000110000001111 ;
ROM[494] <=  32'b01010001000001100101110000010011 ;
ROM[495] <=  32'b01000000000000000000000000000000 ;
ROM[496] <=  32'b00000000000000000000000000000000 ;
ROM[497] <=  32'b00000001001110010110010001001111 ;
ROM[498] <=  32'b10011001010100000111101101111010 ;
ROM[499] <=  32'b10111101000101000100001100101111 ;
ROM[500] <=  32'b01001011111101010001000111010001 ;
ROM[501] <=  32'b00101111000000010100010001001001 ;
ROM[502] <=  32'b00111001001011010101000100000000 ;
ROM[503] <=  32'b01100111111001111001010000111010 ;
ROM[504] <=  32'b01110000000001100111010100010000 ;
ROM[505] <=  32'b10101001010001001011100101000100 ;
ROM[506] <=  32'b01110110100100101001010001010001 ;
ROM[507] <=  32'b00011111101011011100110110010100 ;
ROM[508] <=  32'b00111101010110100100011000000000 ;
ROM[509] <=  32'b00000000000000000000000000000001 ;
ROM[510] <=  32'b00111001011001000100111110011001 ;
ROM[511] <=  32'b01010000101100001001010011100100 ;
ROM[512] <=  32'b01010100010001100000000110001111 ;
ROM[513] <=  32'b11000101000100100000101111111100 ;
ROM[514] <=  32'b10110101010000111011010111100100 ;
ROM[515] <=  32'b10101000010100001100010101110000 ;
ROM[516] <=  32'b11011101100101000011000101110000 ;
ROM[517] <=  32'b00101110110001010000111001010001 ;
ROM[518] <=  32'b10010100110010010100010001011101 ;
ROM[519] <=  32'b11001010111100000101000100100010 ;
ROM[520] <=  32'b00001010001100100101010001000100 ;
ROM[521] <=  32'b10111101100111111011000000000000 ;
ROM[522] <=  32'b00000000000000000000000100111001 ;
ROM[523] <=  32'b01100100010011111001100101010000 ;
ROM[524] <=  32'b11101101100101101111101010010100 ;
ROM[525] <=  32'b01000111110111110001010011010101 ;
ROM[526] <=  32'b00010010001010111001010001111001 ;
ROM[527] <=  32'b01000010110111101101100000010000 ;
ROM[528] <=  32'b01001111111110101100010000111100 ;
ROM[529] <=  32'b11010100000001111011111011010110 ;
ROM[530] <=  32'b10010101000010001001010001101000 ;
ROM[531] <=  32'b00111101010000111110101010001011 ;
ROM[532] <=  32'b10011110010100010010001011001011 ;
ROM[533] <=  32'b11101011100101000100100001110011 ;
ROM[534] <=  32'b11000000000001010000100010100001 ;
ROM[535] <=  32'b10100101110110000000000000000000 ;
ROM[536] <=  32'b00000000000000000101000011101110 ;
ROM[537] <=  32'b11111100111001101101010001001000 ;
ROM[538] <=  32'b00000100001001100111010100010010 ;
ROM[539] <=  32'b00100011010100100110100101000011 ;
ROM[540] <=  32'b00110100001101110001000100000000 ;
ROM[541] <=  32'b00000000000000000000000000010011 ;
ROM[542] <=  32'b10010110010001001111100110010100 ;
ROM[543] <=  32'b11100101100100010011111001100101 ;
ROM[544] <=  32'b01000011100001010010100001011011 ;
ROM[545] <=  32'b01010001000111100111010101011001 ;
ROM[546] <=  32'b10010100010010001101011000111100 ;
ROM[547] <=  32'b11100101000010100010010010111101 ;
ROM[548] <=  32'b01001100000000000000000000000000 ;
ROM[549] <=  32'b00000000010100001110011001110110 ;
ROM[550] <=  32'b11011010000101000100011111001011 ;
ROM[551] <=  32'b01011000100001010001001000111111 ;
ROM[552] <=  32'b01101101100011010100010000011101 ;
ROM[553] <=  32'b10100001110011110101000001010011 ;
ROM[554] <=  32'b00011101110101011101010000011000 ;
ROM[555] <=  32'b01000101100001100100010100001100 ;
ROM[556] <=  32'b10101010010110011111000101000100 ;
ROM[557] <=  32'b00011010011110101011111001010001 ;
ROM[558] <=  32'b00011111001001001111001000010100 ;
ROM[559] <=  32'b01000110101100001110100111000101 ;
ROM[560] <=  32'b00000101100000110111000011001100 ;
ROM[561] <=  32'b00000000000000000000000000000000 ;
ROM[562] <=  32'b01010000101100101110110001110001 ;
ROM[563] <=  32'b01010100010000011010000100110011 ;
ROM[564] <=  32'b11000101000100011110110101100001 ;
ROM[565] <=  32'b00100001010001000111001100101110 ;
ROM[566] <=  32'b10110101010100010000010000101010 ;
ROM[567] <=  32'b00000001010101000011110110110110 ;
ROM[568] <=  32'b11110110000001010001000000111101 ;
ROM[569] <=  32'b11110100100100010100010001010001 ;
ROM[570] <=  32'b10111010001001110101000100011011 ;
ROM[571] <=  32'b10001001010111111001010000111110 ;
ROM[572] <=  32'b00111111101001001011000000000000 ;
ROM[573] <=  32'b00000000000000000000000100111111 ;
ROM[574] <=  32'b10111000001011001101110101010000 ;
ROM[575] <=  32'b00100110101100101000000001010100 ;
ROM[576] <=  32'b00110110101000011110110111100101 ;
ROM[577] <=  32'b00010001010001100100000010011001 ;
ROM[578] <=  32'b01000100100000100110010101101110 ;
ROM[579] <=  32'b01010001000110011001011110101100 ;
ROM[580] <=  32'b11010100010001001000001111110101 ;
ROM[581] <=  32'b00100101000100001011001111110101 ;
ROM[582] <=  32'b10110001010001000011110111000101 ;
ROM[583] <=  32'b11001111010100010000010010000001 ;
ROM[584] <=  32'b00010100010101000001111110100101 ;
ROM[585] <=  32'b11001001110100000000000000000000 ;
ROM[586] <=  32'b00000000000000010011111111101001 ;
ROM[587] <=  32'b00100100010011100100111001011001 ;
ROM[588] <=  32'b00010011111001100101010000011101 ;
ROM[589] <=  32'b11011101101100101010010100001110 ;
ROM[590] <=  32'b01101011101101011101100101000100 ;
ROM[591] <=  32'b00101011100011110110100101010001 ;
ROM[592] <=  32'b00001111000101111001010111010100 ;
ROM[593] <=  32'b01000010101101110100100111010101 ;
ROM[594] <=  32'b00010000001011111011010000111001 ;
ROM[595] <=  32'b01000011110000001110100100000000 ;
ROM[596] <=  32'b01010000110011011111000110110000 ;
ROM[597] <=  32'b11010100000110110010001000011100 ;
ROM[598] <=  32'b11010101000001010011111011011000 ;
ROM[599] <=  32'b10111001001110010110010001001111 ;
ROM[600] <=  32'b10011001010011100101100100010011 ;
ROM[601] <=  32'b11100110010100111001011001000100 ;
ROM[602] <=  32'b11111001100101010000100111111100 ;
ROM[603] <=  32'b11010010110010010100001101010111 ;
ROM[604] <=  32'b00111010010111100101000011110000 ;
ROM[605] <=  32'b10111110101001100101010000111100 ;
ROM[606] <=  32'b11111000011100010010010100001110 ;
ROM[607] <=  32'b10000111110000011101010101000011 ;
ROM[608] <=  32'b01011101010000110010111001010000 ;
ROM[609] <=  32'b10101101010011001101010101010100 ;
ROM[610] <=  32'b00011100111100111111001111000100 ;
ROM[611] <=  32'b11100101100100010011111001100101 ;
ROM[612] <=  32'b00111001011001000100111110011001 ;
*/

end

always @(posedge clk)
begin
out=ROM[addr];
end
endmodule




module COUNTER_LAYER_1024_cycles (clk, count_temp);
input clk;
output reg [9:0] count_temp;
initial begin count_temp <=10'b0000000000; end
always @ (posedge clk)
begin 
count_temp <= count_temp +10'b0000000001;
end
endmodule




module WrapperForFPGA(clk,AXIoutput );

input clk;
output [31:0] AXIoutput;

wire [9:0] addr;
wire [31:0] AXIinput;

COUNTER_LAYER_1024_cycles CounterInstance (clk, addr);
ROM_FPGA_Input  ROMInstance (AXIinput, addr, clk);
happy   happyInstance (clk,  AXIinput, AXIoutput);

endmodule



module WrapperForFPGA_TB();

reg clk ;
wire [31:0] AXIoutput;

WrapperForFPGA  wrapperInstance (clk,AXIoutput );

always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
endmodule
