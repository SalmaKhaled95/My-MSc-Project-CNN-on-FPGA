//line1 bla.v
module TB_bla();

reg clk;
reg rst_Controller;

reg [33:0] DataIn0 , DataIn1 , DataIn2 , DataIn3 ;
localparam period = 100; 
wire [3:0] FinalAnswer;
happy  otta (clk, rst_Controller,FinalAnswer,  DataIn0 , DataIn1 , DataIn2 , DataIn3);
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end
initial 
        begin
		
	    rst_Controller = 1;
		#20;
		rst_Controller = 0;
		
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0101000001100100000000000000000000;
DataIn3   <=34'b0101000001111100000000000000000000;
#period;
DataIn0   <=34'b0101000011000010010000000000000000;
DataIn1   <=34'b0101000011000010010000000000000000;
DataIn2   <=34'b0101000011010000000000000000000000;
DataIn3   <=34'b0101000010101011000000000000000000;
#period;
DataIn0   <=34'b0101000010100100000000000000000000;
DataIn1   <=34'b0100111111100000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0101000001010100000000000000000000;
DataIn1   <=34'b0101000010101011000000000000000000;
DataIn2   <=34'b0101000011011110100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011010110010000000000000000;
#period;
DataIn0   <=34'b0101000011011101100000000000000000;
DataIn1   <=34'b0101000011000101110000000000000000;
DataIn2   <=34'b0101000010000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0101000001100000000000000000000000;
#period;
DataIn0   <=34'b0101000011001100110000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011001110000000000000000;
DataIn3   <=34'b0101000010010110000000000000000000;
#period;
DataIn0   <=34'b0101000001011100000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0101000010100100000000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000010110100000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0101000010011101000000000000000000;
DataIn3   <=34'b0101000011001111110000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000010110110100000000000000000;
DataIn2   <=34'b0101000010101001100000000000000000;
DataIn3   <=34'b0101000011010001110000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011100110000000000000000;
DataIn1   <=34'b0101000010101010100000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0101000011001011000000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011010010100000000000000000;
DataIn3   <=34'b0101000011000100110000000000000000;
#period;
DataIn0   <=34'b0101000011000100110000000000000000;
DataIn1   <=34'b0101000010001101000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0101000001001100000000000000000000;
#period;
DataIn0   <=34'b0101000001111010000000000000000000;
DataIn1   <=34'b0101000011010010000000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011001010110000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0100111111100000000000000000000000;
DataIn2   <=34'b0101000011001011100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000010101100100000000000000000;
DataIn2   <=34'b0101000010100001100000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0101000011000000000000000000000000;
DataIn2   <=34'b0101000011011111000000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011010101000000000000000000;
DataIn2   <=34'b0101000010100110000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0101000010001111000000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000001111010000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0101000010101001100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011000110010000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0101000010101000000000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011100000000000000000000;
DataIn1   <=34'b0101000001110000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0101000001110010000000000000000000;
DataIn3   <=34'b0101000011011100000000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011000110010000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0101000010100000000000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011001110100000000000000000;
DataIn1   <=34'b0101000000111000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0101000011001001100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011000000000000000000000;
DataIn3   <=34'b0101000001010000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0101000001011000000000000000000000;
DataIn1   <=34'b0101000011011010000000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000001111010000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0101000010100101100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000001100010000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0101000001100100000000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000001111010000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0101000010010000000000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000001100010000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0101000000000000000000000000000000;
DataIn1   <=34'b0101000011001000110000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000001111010000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0101000010010000000000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000001100010000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0101000010101111000000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011010010000000000000000000;
DataIn2   <=34'b0101000001010000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0101000001100000000000000000000000;
DataIn3   <=34'b0101000011010100010000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011000101100000000000000000;
DataIn3   <=34'b0100111111100000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0101000001011100000000000000000000;
DataIn2   <=34'b0101000011010011100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011010010100000000000000000;
DataIn3   <=34'b0101000010100001000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0101000001101010000000000000000000;
DataIn2   <=34'b0101000011001000010000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011101010000000000000000;
DataIn2   <=34'b0101000001111110000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0101000010011100000000000000000000;
DataIn3   <=34'b0101000011010101000000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011010000100000000000000000;
#period;
DataIn0   <=34'b0101000010010000000000000000000000;
DataIn1   <=34'b0101000010010000000000000000000000;
DataIn2   <=34'b0101000010000010000000000000000000;
DataIn3   <=34'b0101000010001001000000000000000000;
#period;
DataIn0   <=34'b0101000010010000000000000000000000;
DataIn1   <=34'b0101000011010100010000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011001010110000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0101000010101011000000000000000000;
#period;
DataIn0   <=34'b0101000011011100110000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011010010000000000000000;
DataIn3   <=34'b0101000011011100110000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000010101011000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0101000010111001000000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011011110000000000000000;
#period;
DataIn0   <=34'b0101000010101011000000000000000000;
DataIn1   <=34'b0101000001001100000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0101000001010100000000000000000000;
DataIn1   <=34'b0101000011001101100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111100000000000000000;
DataIn2   <=34'b0101000011011100110000000000000000;
DataIn3   <=34'b0101000010100011000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0101000001000000000000000000000000;
DataIn2   <=34'b0101000010100110000000000000000000;
DataIn3   <=34'b0101000011000100100000000000000000;
#period;
DataIn0   <=34'b0101000011011111100000000000000000;
DataIn1   <=34'b0101000011011111110000000000000000;
DataIn2   <=34'b0101000011011111100000000000000000;
DataIn3   <=34'b0101000011011111110000000000000000;
#period;
DataIn0   <=34'b0101000011000100100000000000000000;
DataIn1   <=34'b0101000001100110000000000000000000;
DataIn2   <=34'b0101000001011100000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;
DataIn0   <=34'b0000000000000000000000000000000000;
DataIn1   <=34'b0000000000000000000000000000000000;
DataIn2   <=34'b0000000000000000000000000000000000;
DataIn3   <=34'b0000000000000000000000000000000000;
#period;

		
		        end
				endmodule


