module MAC_9 (A, B, clk, Z, MAC_start, MAC_end, resetTheCounter);
input [65:0] A;
input [65:0] B;
output  [65:0] Z;
input clk;
input MAC_start, MAC_end;
wire [65:0] R;
input resetTheCounter;
DoublePointMultiplier MultiplierInstance (clk, A , B , R );	
AdderAcc_9 AdderAcc9 (R, clk, Z, MAC_start, MAC_end, resetTheCounter);

endmodule


module AdderAcc_9 (A, clk, Z, MAC_start, MAC_end, resetTheCounter);
input [65:0] A;
input clk;
input MAC_start, MAC_end;
output [65:0] Z;
reg [65:0] R1;
wire [65:0] TempOut;
reg [65:0] Acc = 66'b0;
wire [7:0] count_temp;
wire startCounter, endCounter;
assign startCounter = (MAC_start && !MAC_end)? 1'b1: 1'b0;
input resetTheCounter;
COUNTER_LAYER_222_cycles TheCounter (clk, resetTheCounter, count_temp, startCounter,endCounter);
DoubleAdder AdderInstance (clk,  R1 ,  Acc ,  TempOut  ); 

always @ (posedge clk)
begin 

if (count_temp ==  13  ) begin   Acc = TempOut; /*$display(",  1 , TempOut = %b", TempOut); */ end
else if (count_temp ==  26  ) begin   Acc = TempOut; /*$display(",  2 , TempOut = %b", TempOut); */ end
else if (count_temp ==  39  ) begin   Acc = TempOut; /*$display(",  3 , TempOut = %b", TempOut); */ end
else if (count_temp ==  52  ) begin   Acc = TempOut; /*$display(",  4 , TempOut = %b", TempOut); */ end
else if (count_temp ==  65  ) begin   Acc = TempOut; /*$display(",  5 , TempOut = %b", TempOut); */ end
else if (count_temp ==  78  ) begin   Acc = TempOut; /*$display(",  6 , TempOut = %b", TempOut); */ end
else if (count_temp ==  91  ) begin   Acc = TempOut; /*$display(",  7 , TempOut = %b", TempOut); */ end
else if (count_temp ==  104  ) begin   Acc = TempOut; /*$display(",  8 , TempOut = %b", TempOut); */ end
//if (count_temp ==  117  ) begin   Acc = TempOut; /*$display(",  9 , TempOut = %b", TempOut); */ end
if (!MAC_start && !MAC_end ) begin Acc = 0; end
R1= A; 
end 

assign Z = (MAC_end)? TempOut: 66'bz;
endmodule



module AdderAcc_5 (A, clk, Z, MAC_start, MAC_end, resetTheCounter);
input [65:0] A;
input clk;
input MAC_start, MAC_end;
output [65:0] Z;
reg [65:0] R1;
wire [65:0] TempOut;
reg [65:0] Acc = 66'b0;
wire [6:0] count_temp;
wire startCounter, endCounter;
assign startCounter = (MAC_start && !MAC_end)? 1'b1: 1'b0;
input resetTheCounter;
COUNTER_LAYER_65_cycles TheCounter (clk,resetTheCounter, count_temp, startCounter,endCounter); //66 cycles
DoubleAdder AdderInstance (clk,  R1 ,  Acc ,  TempOut  );

always @ (posedge clk)
begin 

if (resetTheCounter) begin Acc = 0; end
else if (count_temp ==  13  ) begin   Acc = TempOut; /*$display(",  1 , TempOut = %b", TempOut); */ end
else if (count_temp ==  26  ) begin   Acc = TempOut; /*$display(",  2 , TempOut = %b", TempOut); */ end
else if (count_temp ==  39  ) begin   Acc = TempOut; /*$display(",  3 , TempOut = %b", TempOut); */ end
else if (count_temp ==  52  ) begin   Acc = TempOut; /*$display(",  4 , TempOut = %b", TempOut); */ end
else if (count_temp ==  65  ) begin   Acc = TempOut; /*$display(",  5 , TempOut = %b", TempOut); */ end
else if (!MAC_start && !MAC_end ) begin Acc = 0; end
R1= A; 
end 

assign Z = (MAC_end)? TempOut: 66'bz;
endmodule



/*
module COUNTER_LAYER_5550_cycles(clk, count_temp, startOfLayer,endofLayer, bigaddress222);
input clk;
input startOfLayer;
output reg [4:0] bigaddress222;
output endofLayer;
output reg [12:0] count_temp;
initial begin count_temp <=13'b0000000000000; end
always @ (posedge clk)
begin 
if(startOfLayer) begin count_temp <= count_temp +13'b0000000000001; end
//1010110101110 --> 2**12 + 2**10 + 2**8 + 2**7 + 2 **5 + 2**3 + 2**2 + 2**1
end
assign endofLayer = ((((!count_temp[0] && count_temp[1] )&& (count_temp[2] && count_temp[3])) && 
((!count_temp[4] && count_temp[5] )&& (!count_temp[6] && count_temp[7] )))&& 
(((count_temp[8] && !count_temp[9] )&& (count_temp[10] && !count_temp[11] ))&& 
count_temp[12] )) ;


always @ (posedge clk)
begin 
if (count_temp == 0) begin bigaddress222 <= 1; end
else if (count_temp == 222) begin bigaddress222 <= 2 ; end 
else if (count_temp == 444) begin bigaddress222 <= 3 ; end 
else if (count_temp == 666) begin bigaddress222 <= 4 ; end 
else if (count_temp == 888) begin bigaddress222 <= 5 ; end 
else if (count_temp == 1110) begin bigaddress222 <= 6 ; end 
else if (count_temp == 1332) begin bigaddress222 <= 7 ; end 
else if (count_temp == 1554) begin bigaddress222 <= 8 ; end 
else if (count_temp == 1776) begin bigaddress222 <= 9 ; end 
else if (count_temp == 1998) begin bigaddress222 <= 10 ; end 
else if (count_temp == 2220) begin bigaddress222 <= 11 ; end 
else if (count_temp == 2442) begin bigaddress222 <= 12 ; end 
else if (count_temp == 2664) begin bigaddress222 <= 13 ; end 
else if (count_temp == 2886) begin bigaddress222 <= 14 ; end 
else if (count_temp == 3108) begin bigaddress222 <= 15 ; end 
else if (count_temp == 3330) begin bigaddress222 <= 16 ; end 
else if (count_temp == 3552) begin bigaddress222 <= 17 ; end 
else if (count_temp == 3774) begin bigaddress222 <= 18 ; end 
else if (count_temp == 3996) begin bigaddress222 <= 19 ; end 
else if (count_temp == 4218) begin bigaddress222 <= 20 ; end 
else if (count_temp == 4440) begin bigaddress222 <= 21 ; end 
else if (count_temp == 4662) begin bigaddress222 <= 22 ; end 
else if (count_temp == 4884) begin bigaddress222 <= 23 ; end 
else if (count_temp == 5106) begin bigaddress222 <= 24 ; end 
else if (count_temp == 5328) begin bigaddress222 <= 25 ; end 
end
endmodule

*/

module COUNTER_LAYER_5552_cycles_2(clk, count_temp, startOfLayer,endofLayer, bigaddress222);
input clk;
input startOfLayer;
output reg [4:0] bigaddress222;
output endofLayer;
output reg [12:0] count_temp;
initial begin count_temp <=13'b0000000000000; end
always @ (posedge clk)
begin 
if(startOfLayer) begin count_temp <= count_temp +13'b0000000000001; end
//1010110101110 --> 2**12 + 2**10 + 2**8 + 2**7 + 2 **5 + 2**3 + 2**2 + 2**1
end
assign endofLayer = ((((!count_temp[0] && !count_temp[1] )&& (!count_temp[2] && !count_temp[3])) && 
((count_temp[4] && count_temp[5] )&& (!count_temp[6] && count_temp[7] )))&& 
(((count_temp[8] && !count_temp[9] )&& (count_temp[10] && !count_temp[11] ))&& 
count_temp[12] )) ;
///1010110110000

always @ (posedge clk)
begin 
if (count_temp == 0) begin bigaddress222 <= 1; end
else if (count_temp == 222) begin bigaddress222 <= 2 ; end 
else if (count_temp == 444) begin bigaddress222 <= 3 ; end 
else if (count_temp == 666) begin bigaddress222 <= 4 ; end 
else if (count_temp == 888) begin bigaddress222 <= 5 ; end 
else if (count_temp == 1110) begin bigaddress222 <= 6 ; end 
else if (count_temp == 1332) begin bigaddress222 <= 7 ; end 
else if (count_temp == 1554) begin bigaddress222 <= 8 ; end 
else if (count_temp == 1776) begin bigaddress222 <= 9 ; end 
else if (count_temp == 1998) begin bigaddress222 <= 10 ; end 
else if (count_temp == 2220) begin bigaddress222 <= 11 ; end 
else if (count_temp == 2442) begin bigaddress222 <= 12 ; end 
else if (count_temp == 2664) begin bigaddress222 <= 13 ; end 
else if (count_temp == 2886) begin bigaddress222 <= 14 ; end 
else if (count_temp == 3108) begin bigaddress222 <= 15 ; end 
else if (count_temp == 3330) begin bigaddress222 <= 16 ; end 
else if (count_temp == 3552) begin bigaddress222 <= 17 ; end 
else if (count_temp == 3774) begin bigaddress222 <= 18 ; end 
else if (count_temp == 3996) begin bigaddress222 <= 19 ; end 
else if (count_temp == 4218) begin bigaddress222 <= 20 ; end 
else if (count_temp == 4440) begin bigaddress222 <= 21 ; end 
else if (count_temp == 4662) begin bigaddress222 <= 22 ; end 
else if (count_temp == 4884) begin bigaddress222 <= 23 ; end 
else if (count_temp == 5106) begin bigaddress222 <= 24 ; end 
else if (count_temp == 5328) begin bigaddress222 <= 25 ; end 
end
endmodule



module COUNTER_LAYER_1112_cycles_2(clk, count_temp, startOfLayer,endofLayer, bigaddress222);
input clk;
input startOfLayer;
output reg [2:0] bigaddress222;
output endofLayer;
output reg [10:0] count_temp;
initial begin count_temp <=11'b00000000000; end
always @ (posedge clk)
begin 
if(startOfLayer) begin count_temp <= count_temp +11'b00000000001; end
end
assign endofLayer = ((((!count_temp[0] && !count_temp[1] )&& (!count_temp[2] && count_temp[3])) && 
((count_temp[4] && !count_temp[5] )&& (count_temp[6] && !count_temp[7] )))&& 
(((!count_temp[8] && !count_temp[9] )&& count_temp[10]))) ;


//10001011000

always @ (posedge clk)
begin 
if (count_temp == 0) begin bigaddress222 <= 1; end
else if (count_temp == 222) begin bigaddress222 <= 2 ; end 
else if (count_temp == 444) begin bigaddress222 <= 3 ; end 
else if (count_temp == 666) begin bigaddress222 <= 4 ; end 
else if (count_temp == 888) begin bigaddress222 <= 5 ; end 
end
endmodule



module COUNTER_LAYER_65_cycles(clk, RST65, count_temp, startOfLayer,endofLayer);
input clk, RST65;
input startOfLayer;
output endofLayer;
output reg [6:0] count_temp;
initial begin count_temp <=7'b0000000; end
always @ (posedge clk)
begin 
if (RST65) begin count_temp <=7'b0000000; end
else if(startOfLayer) begin count_temp <= count_temp +7'b0000001; end
end
assign endofLayer = (((count_temp[0] && !count_temp[1] )&& (!count_temp[2] && !count_temp[3])) && 
((!count_temp[4] && !count_temp[5] )&& (count_temp[6]))) ;
endmodule




module COUNTER_LAYER_200_cycles(clk, RST157, count_temp, startOfLayer,endofLayer);
//2**7 + 2**6 + 2**3
input clk, RST157;
input startOfLayer;
output endofLayer;
output reg [7:0] count_temp;
initial begin count_temp <=8'b00000000; end
always @ (posedge clk)
begin 
if (RST157) begin count_temp <=8'b00000000; end
else if(startOfLayer) begin count_temp <= count_temp +8'b00000001; end
end
assign endofLayer = (((!count_temp[0] && !count_temp[1] )&& (!count_temp[2] && count_temp[3])) && 
((!count_temp[4] && !count_temp[5] )&& (count_temp[6] && count_temp[7]))) ;
endmodule



module COUNTER_LAYER_222_cycles(clk, resetTheCounter, count_temp, startOfLayer,endofLayer);
//2**7 + 2**6 + 2**4 +  2**3 + 2**2 +2**1
input clk, resetTheCounter;
input startOfLayer;
output endofLayer;
output reg [7:0] count_temp;
initial begin count_temp <=8'b00000000; end
always @ (posedge clk)
begin 
if (resetTheCounter) begin count_temp <=8'b00000000; end
else if(startOfLayer) begin count_temp <= count_temp +8'b00000001; end
end
assign endofLayer = (((!count_temp[0] && count_temp[1] )&& (count_temp[2] && count_temp[3])) && 
((count_temp[4] && !count_temp[5] )&& (count_temp[6] && count_temp[7]))) ;
endmodule



/*
module SUPERMUXMODULECONV2( In0 , In1 , In2 , In3 , In4 , In5 , In6 , In7 , In8 , In9 , In10 , In11 , In12 , In13 , In14 , In15 , 
 In16, In17, In18, In19, In20, In21, In22, In23, In24 ,sel,out );

input [65:0] In0 , In1 , In2 , In3 , In4, In5 , In6 , In7 , In8 , In9 , In10 , In11 , In12 , In13 , In14 , In15 ,  In16, In17, In18, In19, In20, In21, In22, In23, In24 ;
input [12:0] sel;
output [65:0] out;
assign out =

(sel>= 0 && sel< 222 ) ? In0 : 
(sel>= 222 && sel< 444 ) ? In1 :
(sel>= 444 && sel< 666 ) ? In2 :
(sel>= 666 && sel< 888 ) ? In3 :
(sel>= 888 && sel< 1110 ) ? In4 :
(sel>= 1110 && sel< 1332 ) ? In5 :
(sel>= 1332 && sel< 1554 ) ? In6 :
(sel>= 1554 && sel< 1776 ) ? In7 :
(sel>= 1776 && sel< 1998 ) ? In8 :
(sel>= 1998 && sel< 2220 ) ? In9 :
(sel>= 2220 && sel< 2442 ) ? In10 :
(sel>= 2442 && sel< 2664 ) ? In11 :
(sel>= 2664 && sel< 2886 ) ? In12 :
(sel>= 2886 && sel< 3108 ) ? In13 :
(sel>= 3108 && sel< 3330 ) ? In14 :
(sel>= 3330 && sel< 3552 ) ? In15 : 
(sel>= 3552 && sel< 3774 ) ? In16 :
(sel>= 3774 && sel< 3996 ) ? In17 :
(sel>= 3996 && sel< 4218 ) ? In18 :
(sel>= 4218 && sel< 4440 ) ? In19 :
(sel>= 4440 && sel< 4662 ) ? In20 :
(sel>= 4662 && sel< 4884 ) ? In21 :
(sel>= 4884 && sel< 5106 ) ? In22 :
(sel>= 5106 && sel< 5328 ) ? In23 :
(sel>= 5328 && sel< 5550 ) ? In24 :
66'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz; 
endmodule
*/

module SUPERMUXMODULECONV2_new( In0 , In1 , In2 , In3 , In4 , In5 , In6 , In7 , In8 , In9 , In10 , In11 , In12 , In13 , In14 , In15 , 
 In16, In17, In18, In19, In20, In21, In22, In23, In24 ,sel,out );

input [65:0] In0 , In1 , In2 , In3 , In4, In5 , In6 , In7 , In8 , In9 , In10 , In11 , In12 , In13 , In14 , In15 ,  In16, In17, In18, In19, In20, In21, In22, In23, In24 ;
input [4:0] sel;
output reg [65:0] out;

always@(*)
begin
if (sel== 1) begin out = In0 ; end 
else if (sel== 2) begin out = In1 ; end 
else if (sel== 3) begin out = In2 ; end 
else if (sel== 4) begin out = In3 ; end 
else if (sel== 5) begin out = In4 ; end 
else if (sel== 6) begin out = In5 ; end 
else if (sel== 7) begin out = In6 ; end 
else if (sel== 8) begin out = In7 ; end 
else if (sel== 9) begin out = In8 ; end 
else if (sel== 10) begin out = In9 ; end 
else if (sel== 11) begin out = In10 ; end 
else if (sel== 12) begin out = In11 ; end 
else if (sel== 13) begin out = In12 ; end 
else if (sel== 14) begin out = In13 ; end 
else if (sel== 15) begin out = In14 ; end 
else if (sel== 16) begin out = In15 ; end 
else if (sel== 17) begin out = In16 ; end 
else if (sel== 18) begin out = In17 ; end 
else if (sel== 19) begin out = In18 ; end 
else if (sel== 20) begin out = In19 ; end 
else if (sel== 21) begin out = In20 ; end 
else if (sel== 22) begin out = In21 ; end 
else if (sel== 23) begin out = In22 ; end 
else if (sel== 24) begin out = In23 ; end 
else if (sel== 25) begin out = In24 ; end 
end 
/* assign out =

(sel>= 0 && sel< 222 ) ? In0 : 
(sel>= 222 && sel< 444 ) ? In1 :
(sel>= 444 && sel< 666 ) ? In2 :
(sel>= 666 && sel< 888 ) ? In3 :
(sel>= 888 && sel< 1110 ) ? In4 :
(sel>= 1110 && sel< 1332 ) ? In5 :
(sel>= 1332 && sel< 1554 ) ? In6 :
(sel>= 1554 && sel< 1776 ) ? In7 :
(sel>= 1776 && sel< 1998 ) ? In8 :
(sel>= 1998 && sel< 2220 ) ? In9 :
(sel>= 2220 && sel< 2442 ) ? In10 :
(sel>= 2442 && sel< 2664 ) ? In11 :
(sel>= 2664 && sel< 2886 ) ? In12 :
(sel>= 2886 && sel< 3108 ) ? In13 :
(sel>= 3108 && sel< 3330 ) ? In14 :
(sel>= 3330 && sel< 3552 ) ? In15 : 
(sel>= 3552 && sel< 3774 ) ? In16 :
(sel>= 3774 && sel< 3996 ) ? In17 :
(sel>= 3996 && sel< 4218 ) ? In18 :
(sel>= 4218 && sel< 4440 ) ? In19 :
(sel>= 4440 && sel< 4662 ) ? In20 :
(sel>= 4662 && sel< 4884 ) ? In21 :
(sel>= 4884 && sel< 5106 ) ? In22 :
(sel>= 5106 && sel< 5328 ) ? In23 :
(sel>= 5328 && sel< 5550 ) ? In24 :
66'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;  */
endmodule



module SUPERMUXMODULECONV2_new_1_3(  In20, In21, In22, In23, In24 ,sel,out );

input [65:0] In20, In21, In22, In23, In24 ;
input [2:0] sel;
output reg [65:0] out;

always@(*)
begin
if (sel== 1) begin out = In20 ; end 
else if (sel== 2) begin out = In21 ; end 
else if (sel== 3) begin out = In22 ; end 
else if (sel== 4) begin out = In23 ; end 
else if (sel== 5) begin out = In24 ; end 
end 

endmodule




/*
module CONV2LAYER_bla3 (clk, Conv2LayerStart, LayerFinishStage2
,REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143 
, LastRamOutF1_0,LastRamOutF1_1,LastRamOutF1_2,LastRamOutF1_3,LastRamOutF1_4,LastRamOutF1_5,LastRamOutF1_6,LastRamOutF1_7,LastRamOutF1_8,LastRamOutF1_9,LastRamOutF1_10,LastRamOutF1_11,LastRamOutF1_12,LastRamOutF1_13,LastRamOutF1_14,LastRamOutF1_15,LastRamOutF1_16,LastRamOutF1_17,LastRamOutF1_18,LastRamOutF1_19,LastRamOutF1_20,LastRamOutF1_21,LastRamOutF1_22,LastRamOutF1_23,LastRamOutF1_24,LastRamOutF1_25,LastRamOutF1_26,LastRamOutF1_27,LastRamOutF1_28,LastRamOutF1_29,LastRamOutF1_30,LastRamOutF1_31,LastRamOutF1_32,LastRamOutF1_33,LastRamOutF1_34,LastRamOutF1_35,LastRamOutF1_36,LastRamOutF1_37,LastRamOutF1_38,LastRamOutF1_39,LastRamOutF1_40,LastRamOutF1_41,LastRamOutF1_42,LastRamOutF1_43,LastRamOutF1_44,LastRamOutF1_45,LastRamOutF1_46,LastRamOutF1_47,LastRamOutF1_48,LastRamOutF1_49,LastRamOutF1_50,LastRamOutF1_51,LastRamOutF1_52,LastRamOutF1_53,LastRamOutF1_54,LastRamOutF1_55,LastRamOutF1_56,LastRamOutF1_57,LastRamOutF1_58,LastRamOutF1_59,LastRamOutF1_60,LastRamOutF1_61,LastRamOutF1_62,LastRamOutF1_63,LastRamOutF1_64,LastRamOutF1_65,LastRamOutF1_66,LastRamOutF1_67,LastRamOutF1_68,LastRamOutF1_69,LastRamOutF1_70,LastRamOutF1_71,LastRamOutF1_72,LastRamOutF1_73,LastRamOutF1_74,LastRamOutF1_75,LastRamOutF1_76,LastRamOutF1_77,LastRamOutF1_78,LastRamOutF1_79,LastRamOutF1_80,LastRamOutF1_81,LastRamOutF1_82,LastRamOutF1_83,LastRamOutF1_84,LastRamOutF1_85,LastRamOutF1_86,LastRamOutF1_87,LastRamOutF1_88,LastRamOutF1_89,LastRamOutF1_90,LastRamOutF1_91,LastRamOutF1_92,LastRamOutF1_93,LastRamOutF1_94,LastRamOutF1_95,LastRamOutF1_96,LastRamOutF1_97,LastRamOutF1_98,LastRamOutF1_99
, LastRamOutF2_0,LastRamOutF2_1,LastRamOutF2_2,LastRamOutF2_3,LastRamOutF2_4,LastRamOutF2_5,LastRamOutF2_6,LastRamOutF2_7,LastRamOutF2_8,LastRamOutF2_9,LastRamOutF2_10,LastRamOutF2_11,LastRamOutF2_12,LastRamOutF2_13,LastRamOutF2_14,LastRamOutF2_15,LastRamOutF2_16,LastRamOutF2_17,LastRamOutF2_18,LastRamOutF2_19,LastRamOutF2_20,LastRamOutF2_21,LastRamOutF2_22,LastRamOutF2_23,LastRamOutF2_24,LastRamOutF2_25,LastRamOutF2_26,LastRamOutF2_27,LastRamOutF2_28,LastRamOutF2_29,LastRamOutF2_30,LastRamOutF2_31,LastRamOutF2_32,LastRamOutF2_33,LastRamOutF2_34,LastRamOutF2_35,LastRamOutF2_36,LastRamOutF2_37,LastRamOutF2_38,LastRamOutF2_39,LastRamOutF2_40,LastRamOutF2_41,LastRamOutF2_42,LastRamOutF2_43,LastRamOutF2_44,LastRamOutF2_45,LastRamOutF2_46,LastRamOutF2_47,LastRamOutF2_48,LastRamOutF2_49,LastRamOutF2_50,LastRamOutF2_51,LastRamOutF2_52,LastRamOutF2_53,LastRamOutF2_54,LastRamOutF2_55,LastRamOutF2_56,LastRamOutF2_57,LastRamOutF2_58,LastRamOutF2_59,LastRamOutF2_60,LastRamOutF2_61,LastRamOutF2_62,LastRamOutF2_63,LastRamOutF2_64,LastRamOutF2_65,LastRamOutF2_66,LastRamOutF2_67,LastRamOutF2_68,LastRamOutF2_69,LastRamOutF2_70,LastRamOutF2_71,LastRamOutF2_72,LastRamOutF2_73,LastRamOutF2_74,LastRamOutF2_75,LastRamOutF2_76,LastRamOutF2_77,LastRamOutF2_78,LastRamOutF2_79,LastRamOutF2_80,LastRamOutF2_81,LastRamOutF2_82,LastRamOutF2_83,LastRamOutF2_84,LastRamOutF2_85,LastRamOutF2_86,LastRamOutF2_87,LastRamOutF2_88,LastRamOutF2_89,LastRamOutF2_90,LastRamOutF2_91,LastRamOutF2_92,LastRamOutF2_93,LastRamOutF2_94,LastRamOutF2_95,LastRamOutF2_96,LastRamOutF2_97,LastRamOutF2_98,LastRamOutF2_99
, LastRamOutF3_0,LastRamOutF3_1,LastRamOutF3_2,LastRamOutF3_3,LastRamOutF3_4,LastRamOutF3_5,LastRamOutF3_6,LastRamOutF3_7,LastRamOutF3_8,LastRamOutF3_9,LastRamOutF3_10,LastRamOutF3_11,LastRamOutF3_12,LastRamOutF3_13,LastRamOutF3_14,LastRamOutF3_15,LastRamOutF3_16,LastRamOutF3_17,LastRamOutF3_18,LastRamOutF3_19,LastRamOutF3_20,LastRamOutF3_21,LastRamOutF3_22,LastRamOutF3_23,LastRamOutF3_24,LastRamOutF3_25,LastRamOutF3_26,LastRamOutF3_27,LastRamOutF3_28,LastRamOutF3_29,LastRamOutF3_30,LastRamOutF3_31,LastRamOutF3_32,LastRamOutF3_33,LastRamOutF3_34,LastRamOutF3_35,LastRamOutF3_36,LastRamOutF3_37,LastRamOutF3_38,LastRamOutF3_39,LastRamOutF3_40,LastRamOutF3_41,LastRamOutF3_42,LastRamOutF3_43,LastRamOutF3_44,LastRamOutF3_45,LastRamOutF3_46,LastRamOutF3_47,LastRamOutF3_48,LastRamOutF3_49,LastRamOutF3_50,LastRamOutF3_51,LastRamOutF3_52,LastRamOutF3_53,LastRamOutF3_54,LastRamOutF3_55,LastRamOutF3_56,LastRamOutF3_57,LastRamOutF3_58,LastRamOutF3_59,LastRamOutF3_60,LastRamOutF3_61,LastRamOutF3_62,LastRamOutF3_63,LastRamOutF3_64,LastRamOutF3_65,LastRamOutF3_66,LastRamOutF3_67,LastRamOutF3_68,LastRamOutF3_69,LastRamOutF3_70,LastRamOutF3_71,LastRamOutF3_72,LastRamOutF3_73,LastRamOutF3_74,LastRamOutF3_75,LastRamOutF3_76,LastRamOutF3_77,LastRamOutF3_78,LastRamOutF3_79,LastRamOutF3_80,LastRamOutF3_81,LastRamOutF3_82,LastRamOutF3_83,LastRamOutF3_84,LastRamOutF3_85,LastRamOutF3_86,LastRamOutF3_87,LastRamOutF3_88,LastRamOutF3_89,LastRamOutF3_90,LastRamOutF3_91,LastRamOutF3_92,LastRamOutF3_93,LastRamOutF3_94,LastRamOutF3_95,LastRamOutF3_96,LastRamOutF3_97,LastRamOutF3_98,LastRamOutF3_99
, LastRamOutF4_0,LastRamOutF4_1,LastRamOutF4_2,LastRamOutF4_3,LastRamOutF4_4,LastRamOutF4_5,LastRamOutF4_6,LastRamOutF4_7,LastRamOutF4_8,LastRamOutF4_9,LastRamOutF4_10,LastRamOutF4_11,LastRamOutF4_12,LastRamOutF4_13,LastRamOutF4_14,LastRamOutF4_15,LastRamOutF4_16,LastRamOutF4_17,LastRamOutF4_18,LastRamOutF4_19,LastRamOutF4_20,LastRamOutF4_21,LastRamOutF4_22,LastRamOutF4_23,LastRamOutF4_24,LastRamOutF4_25,LastRamOutF4_26,LastRamOutF4_27,LastRamOutF4_28,LastRamOutF4_29,LastRamOutF4_30,LastRamOutF4_31,LastRamOutF4_32,LastRamOutF4_33,LastRamOutF4_34,LastRamOutF4_35,LastRamOutF4_36,LastRamOutF4_37,LastRamOutF4_38,LastRamOutF4_39,LastRamOutF4_40,LastRamOutF4_41,LastRamOutF4_42,LastRamOutF4_43,LastRamOutF4_44,LastRamOutF4_45,LastRamOutF4_46,LastRamOutF4_47,LastRamOutF4_48,LastRamOutF4_49,LastRamOutF4_50,LastRamOutF4_51,LastRamOutF4_52,LastRamOutF4_53,LastRamOutF4_54,LastRamOutF4_55,LastRamOutF4_56,LastRamOutF4_57,LastRamOutF4_58,LastRamOutF4_59,LastRamOutF4_60,LastRamOutF4_61,LastRamOutF4_62,LastRamOutF4_63,LastRamOutF4_64,LastRamOutF4_65,LastRamOutF4_66,LastRamOutF4_67,LastRamOutF4_68,LastRamOutF4_69,LastRamOutF4_70,LastRamOutF4_71,LastRamOutF4_72,LastRamOutF4_73,LastRamOutF4_74,LastRamOutF4_75,LastRamOutF4_76,LastRamOutF4_77,LastRamOutF4_78,LastRamOutF4_79,LastRamOutF4_80,LastRamOutF4_81,LastRamOutF4_82,LastRamOutF4_83,LastRamOutF4_84,LastRamOutF4_85,LastRamOutF4_86,LastRamOutF4_87,LastRamOutF4_88,LastRamOutF4_89,LastRamOutF4_90,LastRamOutF4_91,LastRamOutF4_92,LastRamOutF4_93,LastRamOutF4_94,LastRamOutF4_95,LastRamOutF4_96,LastRamOutF4_97,LastRamOutF4_98,LastRamOutF4_99 
 );

input clk;
input wire [65:0]  REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143; 
input wire [65:0]  REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143; 
input wire [65:0]  REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143; 
input wire [65:0]  REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143; 
input Conv2LayerStart;
output LayerFinishStage2;
wire Conv2LayerFinish, LayerStartStage2;
wire tttt;
wire [12:0] bigaddress;
wire [4:0] bigaddress222;
COUNTER_LAYER_5550_cycles count5550 (clk, bigaddress, Conv2LayerStart,LayerFinishStage2, bigaddress222);
wire [65:0] DataIn;
assign DataIn=66'b0;
output wire [65:0] LastRamOutF1_0,LastRamOutF1_1,LastRamOutF1_2,LastRamOutF1_3,LastRamOutF1_4,LastRamOutF1_5,LastRamOutF1_6,LastRamOutF1_7,LastRamOutF1_8,LastRamOutF1_9,LastRamOutF1_10,LastRamOutF1_11,LastRamOutF1_12,LastRamOutF1_13,LastRamOutF1_14,LastRamOutF1_15,LastRamOutF1_16,LastRamOutF1_17,LastRamOutF1_18,LastRamOutF1_19,LastRamOutF1_20,LastRamOutF1_21,LastRamOutF1_22,LastRamOutF1_23,LastRamOutF1_24,LastRamOutF1_25,LastRamOutF1_26,LastRamOutF1_27,LastRamOutF1_28,LastRamOutF1_29,LastRamOutF1_30,LastRamOutF1_31,LastRamOutF1_32,LastRamOutF1_33,LastRamOutF1_34,LastRamOutF1_35,LastRamOutF1_36,LastRamOutF1_37,LastRamOutF1_38,LastRamOutF1_39,LastRamOutF1_40,LastRamOutF1_41,LastRamOutF1_42,LastRamOutF1_43,LastRamOutF1_44,LastRamOutF1_45,LastRamOutF1_46,LastRamOutF1_47,LastRamOutF1_48,LastRamOutF1_49,LastRamOutF1_50,LastRamOutF1_51,LastRamOutF1_52,LastRamOutF1_53,LastRamOutF1_54,LastRamOutF1_55,LastRamOutF1_56,LastRamOutF1_57,LastRamOutF1_58,LastRamOutF1_59,LastRamOutF1_60,LastRamOutF1_61,LastRamOutF1_62,LastRamOutF1_63,LastRamOutF1_64,LastRamOutF1_65,LastRamOutF1_66,LastRamOutF1_67,LastRamOutF1_68,LastRamOutF1_69,LastRamOutF1_70,LastRamOutF1_71,LastRamOutF1_72,LastRamOutF1_73,LastRamOutF1_74,LastRamOutF1_75,LastRamOutF1_76,LastRamOutF1_77,LastRamOutF1_78,LastRamOutF1_79,LastRamOutF1_80,LastRamOutF1_81,LastRamOutF1_82,LastRamOutF1_83,LastRamOutF1_84,LastRamOutF1_85,LastRamOutF1_86,LastRamOutF1_87,LastRamOutF1_88,LastRamOutF1_89,LastRamOutF1_90,LastRamOutF1_91,LastRamOutF1_92,LastRamOutF1_93,LastRamOutF1_94,LastRamOutF1_95,LastRamOutF1_96,LastRamOutF1_97,LastRamOutF1_98,LastRamOutF1_99; 
output wire [65:0] LastRamOutF2_0,LastRamOutF2_1,LastRamOutF2_2,LastRamOutF2_3,LastRamOutF2_4,LastRamOutF2_5,LastRamOutF2_6,LastRamOutF2_7,LastRamOutF2_8,LastRamOutF2_9,LastRamOutF2_10,LastRamOutF2_11,LastRamOutF2_12,LastRamOutF2_13,LastRamOutF2_14,LastRamOutF2_15,LastRamOutF2_16,LastRamOutF2_17,LastRamOutF2_18,LastRamOutF2_19,LastRamOutF2_20,LastRamOutF2_21,LastRamOutF2_22,LastRamOutF2_23,LastRamOutF2_24,LastRamOutF2_25,LastRamOutF2_26,LastRamOutF2_27,LastRamOutF2_28,LastRamOutF2_29,LastRamOutF2_30,LastRamOutF2_31,LastRamOutF2_32,LastRamOutF2_33,LastRamOutF2_34,LastRamOutF2_35,LastRamOutF2_36,LastRamOutF2_37,LastRamOutF2_38,LastRamOutF2_39,LastRamOutF2_40,LastRamOutF2_41,LastRamOutF2_42,LastRamOutF2_43,LastRamOutF2_44,LastRamOutF2_45,LastRamOutF2_46,LastRamOutF2_47,LastRamOutF2_48,LastRamOutF2_49,LastRamOutF2_50,LastRamOutF2_51,LastRamOutF2_52,LastRamOutF2_53,LastRamOutF2_54,LastRamOutF2_55,LastRamOutF2_56,LastRamOutF2_57,LastRamOutF2_58,LastRamOutF2_59,LastRamOutF2_60,LastRamOutF2_61,LastRamOutF2_62,LastRamOutF2_63,LastRamOutF2_64,LastRamOutF2_65,LastRamOutF2_66,LastRamOutF2_67,LastRamOutF2_68,LastRamOutF2_69,LastRamOutF2_70,LastRamOutF2_71,LastRamOutF2_72,LastRamOutF2_73,LastRamOutF2_74,LastRamOutF2_75,LastRamOutF2_76,LastRamOutF2_77,LastRamOutF2_78,LastRamOutF2_79,LastRamOutF2_80,LastRamOutF2_81,LastRamOutF2_82,LastRamOutF2_83,LastRamOutF2_84,LastRamOutF2_85,LastRamOutF2_86,LastRamOutF2_87,LastRamOutF2_88,LastRamOutF2_89,LastRamOutF2_90,LastRamOutF2_91,LastRamOutF2_92,LastRamOutF2_93,LastRamOutF2_94,LastRamOutF2_95,LastRamOutF2_96,LastRamOutF2_97,LastRamOutF2_98,LastRamOutF2_99; 
output wire [65:0] LastRamOutF3_0,LastRamOutF3_1,LastRamOutF3_2,LastRamOutF3_3,LastRamOutF3_4,LastRamOutF3_5,LastRamOutF3_6,LastRamOutF3_7,LastRamOutF3_8,LastRamOutF3_9,LastRamOutF3_10,LastRamOutF3_11,LastRamOutF3_12,LastRamOutF3_13,LastRamOutF3_14,LastRamOutF3_15,LastRamOutF3_16,LastRamOutF3_17,LastRamOutF3_18,LastRamOutF3_19,LastRamOutF3_20,LastRamOutF3_21,LastRamOutF3_22,LastRamOutF3_23,LastRamOutF3_24,LastRamOutF3_25,LastRamOutF3_26,LastRamOutF3_27,LastRamOutF3_28,LastRamOutF3_29,LastRamOutF3_30,LastRamOutF3_31,LastRamOutF3_32,LastRamOutF3_33,LastRamOutF3_34,LastRamOutF3_35,LastRamOutF3_36,LastRamOutF3_37,LastRamOutF3_38,LastRamOutF3_39,LastRamOutF3_40,LastRamOutF3_41,LastRamOutF3_42,LastRamOutF3_43,LastRamOutF3_44,LastRamOutF3_45,LastRamOutF3_46,LastRamOutF3_47,LastRamOutF3_48,LastRamOutF3_49,LastRamOutF3_50,LastRamOutF3_51,LastRamOutF3_52,LastRamOutF3_53,LastRamOutF3_54,LastRamOutF3_55,LastRamOutF3_56,LastRamOutF3_57,LastRamOutF3_58,LastRamOutF3_59,LastRamOutF3_60,LastRamOutF3_61,LastRamOutF3_62,LastRamOutF3_63,LastRamOutF3_64,LastRamOutF3_65,LastRamOutF3_66,LastRamOutF3_67,LastRamOutF3_68,LastRamOutF3_69,LastRamOutF3_70,LastRamOutF3_71,LastRamOutF3_72,LastRamOutF3_73,LastRamOutF3_74,LastRamOutF3_75,LastRamOutF3_76,LastRamOutF3_77,LastRamOutF3_78,LastRamOutF3_79,LastRamOutF3_80,LastRamOutF3_81,LastRamOutF3_82,LastRamOutF3_83,LastRamOutF3_84,LastRamOutF3_85,LastRamOutF3_86,LastRamOutF3_87,LastRamOutF3_88,LastRamOutF3_89,LastRamOutF3_90,LastRamOutF3_91,LastRamOutF3_92,LastRamOutF3_93,LastRamOutF3_94,LastRamOutF3_95,LastRamOutF3_96,LastRamOutF3_97,LastRamOutF3_98,LastRamOutF3_99; 
output wire [65:0] LastRamOutF4_0,LastRamOutF4_1,LastRamOutF4_2,LastRamOutF4_3,LastRamOutF4_4,LastRamOutF4_5,LastRamOutF4_6,LastRamOutF4_7,LastRamOutF4_8,LastRamOutF4_9,LastRamOutF4_10,LastRamOutF4_11,LastRamOutF4_12,LastRamOutF4_13,LastRamOutF4_14,LastRamOutF4_15,LastRamOutF4_16,LastRamOutF4_17,LastRamOutF4_18,LastRamOutF4_19,LastRamOutF4_20,LastRamOutF4_21,LastRamOutF4_22,LastRamOutF4_23,LastRamOutF4_24,LastRamOutF4_25,LastRamOutF4_26,LastRamOutF4_27,LastRamOutF4_28,LastRamOutF4_29,LastRamOutF4_30,LastRamOutF4_31,LastRamOutF4_32,LastRamOutF4_33,LastRamOutF4_34,LastRamOutF4_35,LastRamOutF4_36,LastRamOutF4_37,LastRamOutF4_38,LastRamOutF4_39,LastRamOutF4_40,LastRamOutF4_41,LastRamOutF4_42,LastRamOutF4_43,LastRamOutF4_44,LastRamOutF4_45,LastRamOutF4_46,LastRamOutF4_47,LastRamOutF4_48,LastRamOutF4_49,LastRamOutF4_50,LastRamOutF4_51,LastRamOutF4_52,LastRamOutF4_53,LastRamOutF4_54,LastRamOutF4_55,LastRamOutF4_56,LastRamOutF4_57,LastRamOutF4_58,LastRamOutF4_59,LastRamOutF4_60,LastRamOutF4_61,LastRamOutF4_62,LastRamOutF4_63,LastRamOutF4_64,LastRamOutF4_65,LastRamOutF4_66,LastRamOutF4_67,LastRamOutF4_68,LastRamOutF4_69,LastRamOutF4_70,LastRamOutF4_71,LastRamOutF4_72,LastRamOutF4_73,LastRamOutF4_74,LastRamOutF4_75,LastRamOutF4_76,LastRamOutF4_77,LastRamOutF4_78,LastRamOutF4_79,LastRamOutF4_80,LastRamOutF4_81,LastRamOutF4_82,LastRamOutF4_83,LastRamOutF4_84,LastRamOutF4_85,LastRamOutF4_86,LastRamOutF4_87,LastRamOutF4_88,LastRamOutF4_89,LastRamOutF4_90,LastRamOutF4_91,LastRamOutF4_92,LastRamOutF4_93,LastRamOutF4_94,LastRamOutF4_95,LastRamOutF4_96,LastRamOutF4_97,LastRamOutF4_98,LastRamOutF4_99; 

///layer300

///////conv2//////



wire xwrite; 
wire xwrite2;
wire  CONV2_MAC_start, CONV2_MAC_end;
wire [7:0] CONV2_counter;
wire [65:0] In1_CONV2_ROMout , In1_CONV2_ROMout1 , In1_CONV2_ROMout2, In1_CONV2_ROMout3;

wire [3:0] CONV2_address; 
wire [65:0] In1_CONV2_MUXout0,In1_CONV2_MUXout1, In1_CONV2_MUXout10,In1_CONV2_MUXout11;
wire [65:0] In1_CONV2_MACoutF1_0,In1_CONV2_MACoutF1_1,In1_CONV2_MACoutF1_10,In1_CONV2_MACoutF1_11;
wire [65:0] In1_CONV2_MACoutF2_0,In1_CONV2_MACoutF2_1,In1_CONV2_MACoutF2_10,In1_CONV2_MACoutF2_11;
wire [65:0] In1_CONV2_MACoutF3_0,In1_CONV2_MACoutF3_1,In1_CONV2_MACoutF3_10,In1_CONV2_MACoutF3_11;
wire [65:0] In1_CONV2_MACoutF4_0,In1_CONV2_MACoutF4_1,In1_CONV2_MACoutF4_10,In1_CONV2_MACoutF4_11;




wire [65:0] In2_CONV2_ROMout, In2_CONV2_ROMout1 , In2_CONV2_ROMout2, In2_CONV2_ROMout3;
wire [65:0] In2_CONV2_MUXout0,In2_CONV2_MUXout1,In2_CONV2_MUXout10,In2_CONV2_MUXout11;
wire [65:0] In2_CONV2_MACoutF1_0,In2_CONV2_MACoutF1_1,In2_CONV2_MACoutF1_10,In2_CONV2_MACoutF1_11;
wire [65:0] In2_CONV2_MACoutF2_0,In2_CONV2_MACoutF2_1,In2_CONV2_MACoutF2_10,In2_CONV2_MACoutF2_11;
wire [65:0] In2_CONV2_MACoutF3_0,In2_CONV2_MACoutF3_1,In2_CONV2_MACoutF3_10,In2_CONV2_MACoutF3_11;
wire [65:0] In2_CONV2_MACoutF4_0,In2_CONV2_MACoutF4_1,In2_CONV2_MACoutF4_10,In2_CONV2_MACoutF4_11;



wire [65:0] In3_CONV2_ROMout, In3_CONV2_ROMout1 , In3_CONV2_ROMout2, In3_CONV2_ROMout3;
wire [65:0] In3_CONV2_MUXout0,In3_CONV2_MUXout1,In3_CONV2_MUXout10,In3_CONV2_MUXout11;
wire [65:0] In3_CONV2_MACoutF1_0,In3_CONV2_MACoutF1_1,In3_CONV2_MACoutF1_10,In3_CONV2_MACoutF1_11;
wire [65:0] In3_CONV2_MACoutF2_0,In3_CONV2_MACoutF2_1,In3_CONV2_MACoutF2_10,In3_CONV2_MACoutF2_11;
wire [65:0] In3_CONV2_MACoutF3_0,In3_CONV2_MACoutF3_1,In3_CONV2_MACoutF3_10,In3_CONV2_MACoutF3_11;
wire [65:0] In3_CONV2_MACoutF4_0,In3_CONV2_MACoutF4_1,In3_CONV2_MACoutF4_10,In3_CONV2_MACoutF4_11;


wire [65:0] In4_CONV2_ROMout, In4_CONV2_ROMout1 , In4_CONV2_ROMout2, In4_CONV2_ROMout3;
wire [65:0] In4_CONV2_MUXout0,In4_CONV2_MUXout1,In4_CONV2_MUXout10,In4_CONV2_MUXout11;

wire [65:0] In4_CONV2_MACoutF1_0,In4_CONV2_MACoutF1_1,In4_CONV2_MACoutF1_10,In4_CONV2_MACoutF1_11;
wire [65:0] In4_CONV2_MACoutF2_0,In4_CONV2_MACoutF2_1,In4_CONV2_MACoutF2_10,In4_CONV2_MACoutF2_11;
wire [65:0] In4_CONV2_MACoutF3_0,In4_CONV2_MACoutF3_1,In4_CONV2_MACoutF3_10,In4_CONV2_MACoutF3_11;
wire [65:0] In4_CONV2_MACoutF4_0,In4_CONV2_MACoutF4_1,In4_CONV2_MACoutF4_10,In4_CONV2_MACoutF4_11;


wire [65:0] Super_1_1_1_1_ch1 , Super_1_2_1_1_ch1 , Super_1_3_1_1_ch1 , Super_2_1_1_1_ch1 , Super_2_2_1_1_ch1 , Super_2_3_1_1_ch1 , Super_3_1_1_1_ch1 , Super_3_2_1_1_ch1 , Super_3_3_1_1_ch1 ;
wire [65:0] Super_1_1_1_2_ch1 , Super_1_2_1_2_ch1 , Super_1_3_1_2_ch1 , Super_2_1_1_2_ch1 , Super_2_2_1_2_ch1 , Super_2_3_1_2_ch1 , Super_3_1_1_2_ch1 , Super_3_2_1_2_ch1 , Super_3_3_1_2_ch1 ;
wire [65:0] Super_1_1_2_1_ch1 , Super_1_2_2_1_ch1 , Super_1_3_2_1_ch1 , Super_2_1_2_1_ch1 , Super_2_2_2_1_ch1 , Super_2_3_2_1_ch1 , Super_3_1_2_1_ch1 , Super_3_2_2_1_ch1 , Super_3_3_2_1_ch1 ;
wire [65:0] Super_1_1_2_2_ch1 , Super_1_2_2_2_ch1 , Super_1_3_2_2_ch1 , Super_2_1_2_2_ch1 , Super_2_2_2_2_ch1 , Super_2_3_2_2_ch1 , Super_3_1_2_2_ch1 , Super_3_2_2_2_ch1 , Super_3_3_2_2_ch1 ;


wire [65:0] Super_1_1_1_1_ch2 , Super_1_2_1_1_ch2 , Super_1_3_1_1_ch2 , Super_2_1_1_1_ch2 , Super_2_2_1_1_ch2 , Super_2_3_1_1_ch2 , Super_3_1_1_1_ch2 , Super_3_2_1_1_ch2 , Super_3_3_1_1_ch2  ;
wire [65:0] Super_1_1_1_2_ch2 , Super_1_2_1_2_ch2 , Super_1_3_1_2_ch2 , Super_2_1_1_2_ch2 , Super_2_2_1_2_ch2 , Super_2_3_1_2_ch2 , Super_3_1_1_2_ch2 ,   Super_3_2_1_2_ch2 , Super_3_3_1_2_ch2 ;
wire [65:0] Super_1_1_2_1_ch2 , Super_1_2_2_1_ch2 , Super_1_3_2_1_ch2 , Super_2_1_2_1_ch2 , Super_2_2_2_1_ch2 , Super_2_3_2_1_ch2 , Super_3_1_2_1_ch2 , Super_3_2_2_1_ch2 , Super_3_3_2_1_ch2  ;
wire [65:0] Super_1_1_2_2_ch2 , Super_1_2_2_2_ch2 , Super_1_3_2_2_ch2 , Super_2_1_2_2_ch2 , Super_2_2_2_2_ch2 , Super_2_3_2_2_ch2 , Super_3_1_2_2_ch2 ,  Super_3_2_2_2_ch2 , Super_3_3_2_2_ch2 ;

wire [65:0]  Super_1_1_1_1_ch4 , Super_1_2_1_1_ch4 , Super_1_3_1_1_ch4 , Super_2_1_1_1_ch4 , Super_2_2_1_1_ch4 , Super_2_3_1_1_ch4 , Super_3_1_1_1_ch4 , Super_3_2_1_1_ch4 , Super_3_3_1_1_ch4 ;
wire [65:0]  Super_1_1_1_2_ch4 , Super_1_2_1_2_ch4 , Super_1_3_1_2_ch4 , Super_2_1_1_2_ch4 , Super_2_2_1_2_ch4 , Super_2_3_1_2_ch4 , Super_3_1_1_2_ch4 ,   Super_3_2_1_2_ch4 , Super_3_3_1_2_ch4 ;
wire [65:0]  Super_1_1_2_1_ch4 , Super_1_2_2_1_ch4 , Super_1_3_2_1_ch4 , Super_2_1_2_1_ch4 , Super_2_2_2_1_ch4 , Super_2_3_2_1_ch4 , Super_3_1_2_1_ch4 , Super_3_2_2_1_ch4 , Super_3_3_2_1_ch4 ;
wire [65:0]  Super_1_1_2_2_ch4 , Super_1_2_2_2_ch4 , Super_1_3_2_2_ch4 , Super_2_1_2_2_ch4 , Super_2_2_2_2_ch4 , Super_2_3_2_2_ch4 , Super_3_1_2_2_ch4 ,  Super_3_2_2_2_ch4 , Super_3_3_2_2_ch4  ;


wire [65:0] Super_1_1_1_1_ch3 , Super_1_2_1_1_ch3 , Super_1_3_1_1_ch3 , Super_2_1_1_1_ch3 , Super_2_2_1_1_ch3 , Super_2_3_1_1_ch3 , Super_3_1_1_1_ch3 , Super_3_2_1_1_ch3 , Super_3_3_1_1_ch3 ;
wire [65:0] Super_1_1_1_2_ch3 , Super_1_2_1_2_ch3 , Super_1_3_1_2_ch3 , Super_2_1_1_2_ch3 , Super_2_2_1_2_ch3 , Super_2_3_1_2_ch3 , Super_3_1_1_2_ch3 ,   Super_3_2_1_2_ch3 , Super_3_3_1_2_ch3 ;
wire [65:0] Super_1_1_2_1_ch3 , Super_1_2_2_1_ch3 , Super_1_3_2_1_ch3 , Super_2_1_2_1_ch3 , Super_2_2_2_1_ch3 , Super_2_3_2_1_ch3 , Super_3_1_2_1_ch3 , Super_3_2_2_1_ch3 , Super_3_3_2_1_ch3  ;
wire [65:0] Super_1_1_2_2_ch3 , Super_1_2_2_2_ch3 , Super_1_3_2_2_ch3 , Super_2_1_2_2_ch3 , Super_2_2_2_2_ch3 , Super_2_3_2_2_ch3 , Super_3_1_2_2_ch3 ,  Super_3_2_2_2_ch3 , Super_3_3_2_2_ch3 ;




//wire CONV2_rst;
assign xwrite =1'b0;
assign xwrite2 = Conv2LayerFinish;
assign CONV2_MAC_start = (CONV2_counter >0) ?1'b1 :1'b0;//Conv2LayerStart;
assign CONV2_MAC_end = (CONV2_counter >117) ?1'b1 :1'b0; //117 = 9 * 13
//assign CONV2_rst = (CONV2_counter ==8'b00000000)?1'b1 :1'b0;

wire [65:0] Filter1BIASOUT, Filter2BIASOUT ,Filter3BIASOUT, Filter4BIASOUT;
OneRegister_In1_xBIAS Filter1Bias (clk, xwrite, DataIn, Filter1BIASOUT);
OneRegister_In2_xBIAS Filter2Bias (clk, xwrite, DataIn, Filter2BIASOUT);
OneRegister_In3_xBIAS Filter3Bias (clk, xwrite, DataIn, Filter3BIASOUT);
OneRegister_In4_xBIAS Filter4Bias (clk, xwrite, DataIn, Filter4BIASOUT);


//

reg resetTheCounter;
COUNTER_LAYER_200_cycles Conv2Counter200 (clk, resetTheCounter, CONV2_counter, Conv2LayerStart,bbb);
assign Conv2LayerFinish = (CONV2_counter ==157) ?1'b1 :1'b0;

//channel 1 of all filters


In1_ROM_9x66bit_0 In1_Conv2FilterWeights (clk, CONV2_counter, In1_CONV2_ROMout);
In1_ROM_9x66bit_1 In1_Conv2FilterWeights1 (clk, CONV2_counter, In1_CONV2_ROMout1);
In1_ROM_9x66bit_2 In1_Conv2FilterWeights2 (clk, CONV2_counter, In1_CONV2_ROMout2);
In1_ROM_9x66bit_3 In1_Conv2FilterWeights3 (clk, CONV2_counter, In1_CONV2_ROMout3);


//channel 2 of all filters
In2_ROM_9x66bit_0 In2_Conv2FilterWeights (clk, CONV2_counter, In2_CONV2_ROMout);
In2_ROM_9x66bit_1 In2_Conv2FilterWeights1 (clk, CONV2_counter, In2_CONV2_ROMout1);
In2_ROM_9x66bit_2 In2_Conv2FilterWeights2 (clk, CONV2_counter, In2_CONV2_ROMout2);
In2_ROM_9x66bit_3 In2_Conv2FilterWeights3 (clk, CONV2_counter, In2_CONV2_ROMout3);

//channel 3 of all filters
In3_ROM_9x66bit_0 In3_Conv2FilterWeights (clk, CONV2_counter, In3_CONV2_ROMout);
In3_ROM_9x66bit_1 In3_Conv2FilterWeights1 (clk, CONV2_counter, In3_CONV2_ROMout1);
In3_ROM_9x66bit_2 In3_Conv2FilterWeights2 (clk, CONV2_counter, In3_CONV2_ROMout2);
In3_ROM_9x66bit_3 In3_Conv2FilterWeights3 (clk, CONV2_counter, In3_CONV2_ROMout3);


//channel 4 of all filters
In4_ROM_9x66bit_0 In4_Conv2FilterWeights (clk, CONV2_counter, In4_CONV2_ROMout);
In4_ROM_9x66bit_1 In4_Conv2FilterWeights1 (clk, CONV2_counter, In4_CONV2_ROMout1);
In4_ROM_9x66bit_2 In4_Conv2FilterWeights2 (clk, CONV2_counter, In4_CONV2_ROMout2);
In4_ROM_9x66bit_3 In4_Conv2FilterWeights3 (clk, CONV2_counter, In4_CONV2_ROMout3);

//CONV2_main_fsm Conv2StateMachine (clk, CONV2_rst, CONV2_counter, CONV2_address_0, CONV2_address_1 , CONV2_address_2 , CONV2_address_3 , CONV2_address_4 , CONV2_address_5 , CONV2_address_6 , CONV2_address_7, CONV2_address_8, CONV2_address_9, CONV2_address_10, CONV2_address_11, CONV2_address_12, CONV2_address_13, CONV2_address_14, CONV2_address_15, CONV2_address_16,CONV2_address_17,CONV2_address_18,CONV2_address_19,CONV2_address_20,CONV2_address_21,CONV2_address_22,CONV2_address_23,CONV2_address_24,CONV2_address_25,CONV2_address_26,CONV2_address_27,CONV2_address_28,CONV2_address_29,CONV2_address_30,CONV2_address_31,CONV2_address_32,CONV2_address_33,CONV2_address_34,CONV2_address_35,CONV2_address_36,CONV2_address_37,CONV2_address_38,CONV2_address_39,CONV2_address_40,CONV2_address_41,CONV2_address_42,CONV2_address_43,CONV2_address_44,CONV2_address_45,CONV2_address_46,CONV2_address_47,CONV2_address_48,CONV2_address_49,CONV2_address_50,CONV2_address_51,CONV2_address_52,CONV2_address_53,CONV2_address_54,CONV2_address_55,CONV2_address_56,CONV2_address_57,CONV2_address_58,CONV2_address_59,CONV2_address_60,CONV2_address_61,CONV2_address_62,CONV2_address_63,CONV2_address_64,CONV2_address_65,CONV2_address_66,CONV2_address_67,CONV2_address_68,CONV2_address_69,CONV2_address_70,CONV2_address_71,CONV2_address_72,CONV2_address_73,CONV2_address_74,CONV2_address_75,CONV2_address_76,CONV2_address_77,CONV2_address_78,CONV2_address_79,CONV2_address_80,CONV2_address_81,CONV2_address_82,CONV2_address_83,CONV2_address_84,CONV2_address_85,CONV2_address_86,CONV2_address_87,CONV2_address_88,CONV2_address_89,CONV2_address_90,CONV2_address_91,CONV2_address_92,CONV2_address_93,CONV2_address_94,CONV2_address_95,CONV2_address_96,CONV2_address_97,CONV2_address_98,CONV2_address_99);
CONV2_main_fsm Conv2StateMachine (clk, resetTheCounter, CONV2_counter, CONV2_address);


//0->144 input ,, repeat0->99


//from///

SUPERMUXMODULECONV2_new mux1_1_1_1_ch1 ( REGofMAX1DataOut_F1_0, REGofMAX1DataOut_F1_2 , REGofMAX1DataOut_F1_4 , REGofMAX1DataOut_F1_6 , REGofMAX1DataOut_F1_8 , REGofMAX1DataOut_F1_24 ,
 REGofMAX1DataOut_F1_26 , REGofMAX1DataOut_F1_28 , REGofMAX1DataOut_F1_30 , REGofMAX1DataOut_F1_32 , REGofMAX1DataOut_F1_48 , REGofMAX1DataOut_F1_50 , REGofMAX1DataOut_F1_52 ,
 REGofMAX1DataOut_F1_54, REGofMAX1DataOut_F1_56 , REGofMAX1DataOut_F1_72 , REGofMAX1DataOut_F1_74 , REGofMAX1DataOut_F1_76 , REGofMAX1DataOut_F1_78 , REGofMAX1DataOut_F1_80 ,
 REGofMAX1DataOut_F1_96, REGofMAX1DataOut_F1_98 ,REGofMAX1DataOut_F1_100  , REGofMAX1DataOut_F1_102 , REGofMAX1DataOut_F1_104 , bigaddress222, Super_1_1_1_1_ch1 );
SUPERMUXMODULECONV2_new mux1_2_1_1_ch1 ( REGofMAX1DataOut_F1_1 , REGofMAX1DataOut_F1_3 , REGofMAX1DataOut_F1_5 , REGofMAX1DataOut_F1_7 , REGofMAX1DataOut_F1_9 , REGofMAX1DataOut_F1_25 ,
 REGofMAX1DataOut_F1_27 , REGofMAX1DataOut_F1_29 , REGofMAX1DataOut_F1_31 , REGofMAX1DataOut_F1_33 , REGofMAX1DataOut_F1_49 , REGofMAX1DataOut_F1_51 , REGofMAX1DataOut_F1_53 ,
 REGofMAX1DataOut_F1_55, REGofMAX1DataOut_F1_57 , REGofMAX1DataOut_F1_73 , REGofMAX1DataOut_F1_75 , REGofMAX1DataOut_F1_77 , REGofMAX1DataOut_F1_79 , REGofMAX1DataOut_F1_81 ,
 REGofMAX1DataOut_F1_97, REGofMAX1DataOut_F1_99 , REGofMAX1DataOut_F1_101 , REGofMAX1DataOut_F1_103 ,  REGofMAX1DataOut_F1_105, bigaddress222, Super_1_2_1_1_ch1 );
SUPERMUXMODULECONV2_new mux1_3_1_1_ch1 ( REGofMAX1DataOut_F1_2,  REGofMAX1DataOut_F1_4, REGofMAX1DataOut_F1_6 , REGofMAX1DataOut_F1_8 , REGofMAX1DataOut_F1_10 , REGofMAX1DataOut_F1_26 ,
 REGofMAX1DataOut_F1_28 , REGofMAX1DataOut_F1_30 , REGofMAX1DataOut_F1_32 , REGofMAX1DataOut_F1_34 , REGofMAX1DataOut_F1_50 , REGofMAX1DataOut_F1_52 , REGofMAX1DataOut_F1_54 ,
 REGofMAX1DataOut_F1_56, REGofMAX1DataOut_F1_58 , REGofMAX1DataOut_F1_74 , REGofMAX1DataOut_F1_76 , REGofMAX1DataOut_F1_78 , REGofMAX1DataOut_F1_80 , REGofMAX1DataOut_F1_82 ,
 REGofMAX1DataOut_F1_98, REGofMAX1DataOut_F1_100 , REGofMAX1DataOut_F1_102 , REGofMAX1DataOut_F1_104 , REGofMAX1DataOut_F1_106 , bigaddress222, Super_1_3_1_1_ch1 );
SUPERMUXMODULECONV2_new mux2_1_1_1_ch1 ( REGofMAX1DataOut_F1_12 ,REGofMAX1DataOut_F1_14  , REGofMAX1DataOut_F1_16 , REGofMAX1DataOut_F1_18 , REGofMAX1DataOut_F1_20 , REGofMAX1DataOut_F1_36 ,
 REGofMAX1DataOut_F1_38 , REGofMAX1DataOut_F1_40 , REGofMAX1DataOut_F1_42 , REGofMAX1DataOut_F1_44 , REGofMAX1DataOut_F1_60 , REGofMAX1DataOut_F1_62 , REGofMAX1DataOut_F1_64 ,
 REGofMAX1DataOut_F1_66, REGofMAX1DataOut_F1_68 , REGofMAX1DataOut_F1_84 , REGofMAX1DataOut_F1_86 , REGofMAX1DataOut_F1_88 , REGofMAX1DataOut_F1_90 , REGofMAX1DataOut_F1_92  ,
 REGofMAX1DataOut_F1_108, REGofMAX1DataOut_F1_110 , REGofMAX1DataOut_F1_112 , REGofMAX1DataOut_F1_114 , REGofMAX1DataOut_F1_116 , bigaddress222, Super_2_1_1_1_ch1 );
SUPERMUXMODULECONV2_new mux2_2_1_1_ch1 ( REGofMAX1DataOut_F1_13, REGofMAX1DataOut_F1_15 , REGofMAX1DataOut_F1_17 , REGofMAX1DataOut_F1_19 , REGofMAX1DataOut_F1_21 , REGofMAX1DataOut_F1_37 ,
 REGofMAX1DataOut_F1_39 , REGofMAX1DataOut_F1_41 , REGofMAX1DataOut_F1_43 , REGofMAX1DataOut_F1_45 , REGofMAX1DataOut_F1_61 , REGofMAX1DataOut_F1_63 , REGofMAX1DataOut_F1_65 ,
 REGofMAX1DataOut_F1_67, REGofMAX1DataOut_F1_69 , REGofMAX1DataOut_F1_85 , REGofMAX1DataOut_F1_87 , REGofMAX1DataOut_F1_89 , REGofMAX1DataOut_F1_91 ,REGofMAX1DataOut_F1_93  ,
 REGofMAX1DataOut_F1_109, REGofMAX1DataOut_F1_111 , REGofMAX1DataOut_F1_113 , REGofMAX1DataOut_F1_115 ,REGofMAX1DataOut_F1_117  , bigaddress222, Super_2_2_1_1_ch1 );
SUPERMUXMODULECONV2_new mux2_3_1_1_ch1 ( REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_16  , REGofMAX1DataOut_F1_18 , REGofMAX1DataOut_F1_20 , REGofMAX1DataOut_F1_22 , REGofMAX1DataOut_F1_38 ,
 REGofMAX1DataOut_F1_40 , REGofMAX1DataOut_F1_42 , REGofMAX1DataOut_F1_44 , REGofMAX1DataOut_F1_46 , REGofMAX1DataOut_F1_62 , REGofMAX1DataOut_F1_64 , REGofMAX1DataOut_F1_66 ,
 REGofMAX1DataOut_F1_68, REGofMAX1DataOut_F1_70 , REGofMAX1DataOut_F1_86 , REGofMAX1DataOut_F1_88 , REGofMAX1DataOut_F1_90 , REGofMAX1DataOut_F1_92 , REGofMAX1DataOut_F1_94 ,
 REGofMAX1DataOut_F1_110, REGofMAX1DataOut_F1_112 , REGofMAX1DataOut_F1_114 , REGofMAX1DataOut_F1_116 , REGofMAX1DataOut_F1_118 , bigaddress222, Super_2_3_1_1_ch1 );
SUPERMUXMODULECONV2_new mux3_1_1_1_ch1 ( REGofMAX1DataOut_F1_24, REGofMAX1DataOut_F1_26 , REGofMAX1DataOut_F1_28 , REGofMAX1DataOut_F1_30 , REGofMAX1DataOut_F1_32 , REGofMAX1DataOut_F1_48 ,
 REGofMAX1DataOut_F1_50 , REGofMAX1DataOut_F1_52 , REGofMAX1DataOut_F1_54 , REGofMAX1DataOut_F1_56 , REGofMAX1DataOut_F1_72 , REGofMAX1DataOut_F1_74 , REGofMAX1DataOut_F1_76 ,
 REGofMAX1DataOut_F1_78, REGofMAX1DataOut_F1_80 , REGofMAX1DataOut_F1_96 , REGofMAX1DataOut_F1_98 , REGofMAX1DataOut_F1_100 , REGofMAX1DataOut_F1_102 , REGofMAX1DataOut_F1_104 ,
 REGofMAX1DataOut_F1_120, REGofMAX1DataOut_F1_122 , REGofMAX1DataOut_F1_124 , REGofMAX1DataOut_F1_126 , REGofMAX1DataOut_F1_128 , bigaddress222, Super_3_1_1_1_ch1 );
SUPERMUXMODULECONV2_new mux3_2_1_1_ch1 ( REGofMAX1DataOut_F1_25, REGofMAX1DataOut_F1_27 , REGofMAX1DataOut_F1_29 , REGofMAX1DataOut_F1_31 , REGofMAX1DataOut_F1_33 , REGofMAX1DataOut_F1_49 ,
 REGofMAX1DataOut_F1_51 ,REGofMAX1DataOut_F1_53  , REGofMAX1DataOut_F1_55 , REGofMAX1DataOut_F1_57 , REGofMAX1DataOut_F1_73 , REGofMAX1DataOut_F1_75 , REGofMAX1DataOut_F1_77 ,
REGofMAX1DataOut_F1_79 , REGofMAX1DataOut_F1_81 , REGofMAX1DataOut_F1_97 , REGofMAX1DataOut_F1_99 , REGofMAX1DataOut_F1_101 , REGofMAX1DataOut_F1_103 , REGofMAX1DataOut_F1_105 ,
 REGofMAX1DataOut_F1_121 , REGofMAX1DataOut_F1_123 , REGofMAX1DataOut_F1_125 , REGofMAX1DataOut_F1_127 , REGofMAX1DataOut_F1_129 , bigaddress222, Super_3_2_1_1_ch1 );
SUPERMUXMODULECONV2_new mux3_3_1_1_ch1 ( REGofMAX1DataOut_F1_26, REGofMAX1DataOut_F1_28 , REGofMAX1DataOut_F1_30 , REGofMAX1DataOut_F1_32 , REGofMAX1DataOut_F1_34 , REGofMAX1DataOut_F1_50 ,
REGofMAX1DataOut_F1_52  , REGofMAX1DataOut_F1_54 , REGofMAX1DataOut_F1_56 , REGofMAX1DataOut_F1_58 , REGofMAX1DataOut_F1_74 , REGofMAX1DataOut_F1_76 , REGofMAX1DataOut_F1_78 ,
REGofMAX1DataOut_F1_80 , REGofMAX1DataOut_F1_82 , REGofMAX1DataOut_F1_98 , REGofMAX1DataOut_F1_100 , REGofMAX1DataOut_F1_102 , REGofMAX1DataOut_F1_104 , REGofMAX1DataOut_F1_106 ,
 REGofMAX1DataOut_F1_122 , REGofMAX1DataOut_F1_124 , REGofMAX1DataOut_F1_126 , REGofMAX1DataOut_F1_128 , REGofMAX1DataOut_F1_130 , bigaddress222, Super_3_3_1_1_ch1 );



SUPERMUXMODULECONV2_new mux1_1_1_2_ch1 ( REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_3  , REGofMAX1DataOut_F1_5 , REGofMAX1DataOut_F1_7 , REGofMAX1DataOut_F1_9 , REGofMAX1DataOut_F1_25 ,
REGofMAX1DataOut_F1_27 , REGofMAX1DataOut_F1_29 , REGofMAX1DataOut_F1_31 , REGofMAX1DataOut_F1_33 , REGofMAX1DataOut_F1_49 , REGofMAX1DataOut_F1_51 ,REGofMAX1DataOut_F1_53  ,
 REGofMAX1DataOut_F1_55 ,REGofMAX1DataOut_F1_57  , REGofMAX1DataOut_F1_73 , REGofMAX1DataOut_F1_75 , REGofMAX1DataOut_F1_77 , REGofMAX1DataOut_F1_79 , REGofMAX1DataOut_F1_81 ,
 REGofMAX1DataOut_F1_97, REGofMAX1DataOut_F1_99 , REGofMAX1DataOut_F1_101 , REGofMAX1DataOut_F1_103 , REGofMAX1DataOut_F1_105 , bigaddress222, Super_1_1_1_2_ch1 );
SUPERMUXMODULECONV2_new mux1_2_1_2_ch1 ( REGofMAX1DataOut_F1_2, REGofMAX1DataOut_F1_4 , REGofMAX1DataOut_F1_6 , REGofMAX1DataOut_F1_8 , REGofMAX1DataOut_F1_10 , REGofMAX1DataOut_F1_26 ,
REGofMAX1DataOut_F1_28 , REGofMAX1DataOut_F1_30 , REGofMAX1DataOut_F1_32 , REGofMAX1DataOut_F1_34 , REGofMAX1DataOut_F1_50 , REGofMAX1DataOut_F1_52 ,REGofMAX1DataOut_F1_54  ,
 REGofMAX1DataOut_F1_56 , REGofMAX1DataOut_F1_58 , REGofMAX1DataOut_F1_74 , REGofMAX1DataOut_F1_76 , REGofMAX1DataOut_F1_78 , REGofMAX1DataOut_F1_80 , REGofMAX1DataOut_F1_82 ,
 REGofMAX1DataOut_F1_98, REGofMAX1DataOut_F1_100 , REGofMAX1DataOut_F1_102 , REGofMAX1DataOut_F1_104 , REGofMAX1DataOut_F1_106 , bigaddress222, Super_1_2_1_2_ch1 );
SUPERMUXMODULECONV2_new mux1_3_1_2_ch1 ( REGofMAX1DataOut_F1_3, REGofMAX1DataOut_F1_5 , REGofMAX1DataOut_F1_7 , REGofMAX1DataOut_F1_9 , REGofMAX1DataOut_F1_11 , REGofMAX1DataOut_F1_27 ,
REGofMAX1DataOut_F1_29 , REGofMAX1DataOut_F1_31 , REGofMAX1DataOut_F1_33 , REGofMAX1DataOut_F1_35 , REGofMAX1DataOut_F1_51 , REGofMAX1DataOut_F1_53 , REGofMAX1DataOut_F1_55 ,
 REGofMAX1DataOut_F1_57 , REGofMAX1DataOut_F1_59 , REGofMAX1DataOut_F1_75 , REGofMAX1DataOut_F1_77 , REGofMAX1DataOut_F1_79 , REGofMAX1DataOut_F1_81 , REGofMAX1DataOut_F1_83 ,
 REGofMAX1DataOut_F1_99, REGofMAX1DataOut_F1_101 , REGofMAX1DataOut_F1_103 , REGofMAX1DataOut_F1_105 , REGofMAX1DataOut_F1_107 , bigaddress222, Super_1_3_1_2_ch1 );
SUPERMUXMODULECONV2_new mux2_1_1_2_ch1 ( REGofMAX1DataOut_F1_13, REGofMAX1DataOut_F1_15 , REGofMAX1DataOut_F1_17 , REGofMAX1DataOut_F1_19 , REGofMAX1DataOut_F1_21 , REGofMAX1DataOut_F1_37 ,
REGofMAX1DataOut_F1_39 , REGofMAX1DataOut_F1_41 , REGofMAX1DataOut_F1_43 , REGofMAX1DataOut_F1_45 , REGofMAX1DataOut_F1_61 , REGofMAX1DataOut_F1_63  ,REGofMAX1DataOut_F1_65  ,
 REGofMAX1DataOut_F1_67 , REGofMAX1DataOut_F1_69 , REGofMAX1DataOut_F1_85 , REGofMAX1DataOut_F1_87 , REGofMAX1DataOut_F1_89 , REGofMAX1DataOut_F1_91 , REGofMAX1DataOut_F1_93 ,
 REGofMAX1DataOut_F1_109, REGofMAX1DataOut_F1_111 , REGofMAX1DataOut_F1_113 , REGofMAX1DataOut_F1_115 , REGofMAX1DataOut_F1_117 , bigaddress222, Super_2_1_1_2_ch1 );
SUPERMUXMODULECONV2_new mux2_2_1_2_ch1 ( REGofMAX1DataOut_F1_14, REGofMAX1DataOut_F1_16 , REGofMAX1DataOut_F1_18 , REGofMAX1DataOut_F1_20 , REGofMAX1DataOut_F1_22 , REGofMAX1DataOut_F1_38 ,
REGofMAX1DataOut_F1_40  , REGofMAX1DataOut_F1_42 , REGofMAX1DataOut_F1_44 , REGofMAX1DataOut_F1_46 , REGofMAX1DataOut_F1_62 , REGofMAX1DataOut_F1_64 ,REGofMAX1DataOut_F1_66  ,
 REGofMAX1DataOut_F1_68 , REGofMAX1DataOut_F1_70 , REGofMAX1DataOut_F1_86 , REGofMAX1DataOut_F1_88 , REGofMAX1DataOut_F1_90 , REGofMAX1DataOut_F1_92 , REGofMAX1DataOut_F1_94 ,
 REGofMAX1DataOut_F1_110, REGofMAX1DataOut_F1_112 , REGofMAX1DataOut_F1_114 , REGofMAX1DataOut_F1_116 , REGofMAX1DataOut_F1_118 , bigaddress222, Super_2_2_1_2_ch1 );
SUPERMUXMODULECONV2_new mux2_3_1_2_ch1 ( REGofMAX1DataOut_F1_15, REGofMAX1DataOut_F1_17 , REGofMAX1DataOut_F1_19 , REGofMAX1DataOut_F1_21 , REGofMAX1DataOut_F1_23 , REGofMAX1DataOut_F1_39 ,
REGofMAX1DataOut_F1_41  , REGofMAX1DataOut_F1_43 , REGofMAX1DataOut_F1_45 , REGofMAX1DataOut_F1_47 , REGofMAX1DataOut_F1_63 , REGofMAX1DataOut_F1_65 ,REGofMAX1DataOut_F1_67  ,
 REGofMAX1DataOut_F1_69 , REGofMAX1DataOut_F1_71 , REGofMAX1DataOut_F1_87 , REGofMAX1DataOut_F1_89 , REGofMAX1DataOut_F1_91 , REGofMAX1DataOut_F1_93 , REGofMAX1DataOut_F1_95 ,
 REGofMAX1DataOut_F1_111, REGofMAX1DataOut_F1_113 , REGofMAX1DataOut_F1_115 , REGofMAX1DataOut_F1_117 , REGofMAX1DataOut_F1_119 , bigaddress222, Super_2_3_1_2_ch1 );
SUPERMUXMODULECONV2_new mux3_1_1_2_ch1 ( REGofMAX1DataOut_F1_25, REGofMAX1DataOut_F1_27 , REGofMAX1DataOut_F1_29 , REGofMAX1DataOut_F1_31 , REGofMAX1DataOut_F1_33 , REGofMAX1DataOut_F1_49 ,
REGofMAX1DataOut_F1_51 , REGofMAX1DataOut_F1_53 , REGofMAX1DataOut_F1_55 , REGofMAX1DataOut_F1_57 , REGofMAX1DataOut_F1_73 , REGofMAX1DataOut_F1_75 ,REGofMAX1DataOut_F1_77  ,
 REGofMAX1DataOut_F1_79 , REGofMAX1DataOut_F1_81 , REGofMAX1DataOut_F1_97 , REGofMAX1DataOut_F1_99 , REGofMAX1DataOut_F1_101 , REGofMAX1DataOut_F1_103 , REGofMAX1DataOut_F1_105 ,
REGofMAX1DataOut_F1_121 , REGofMAX1DataOut_F1_123 , REGofMAX1DataOut_F1_125 , REGofMAX1DataOut_F1_127 , REGofMAX1DataOut_F1_129 , bigaddress222, Super_3_1_1_2_ch1 );
SUPERMUXMODULECONV2_new mux3_2_1_2_ch1 ( REGofMAX1DataOut_F1_26, REGofMAX1DataOut_F1_28 , REGofMAX1DataOut_F1_30 , REGofMAX1DataOut_F1_32 , REGofMAX1DataOut_F1_34 , REGofMAX1DataOut_F1_50 ,
REGofMAX1DataOut_F1_52  , REGofMAX1DataOut_F1_54 , REGofMAX1DataOut_F1_56 , REGofMAX1DataOut_F1_58 , REGofMAX1DataOut_F1_74 , REGofMAX1DataOut_F1_76 ,REGofMAX1DataOut_F1_78  ,
 REGofMAX1DataOut_F1_80 , REGofMAX1DataOut_F1_82 , REGofMAX1DataOut_F1_98 , REGofMAX1DataOut_F1_100 , REGofMAX1DataOut_F1_102 , REGofMAX1DataOut_F1_104 ,REGofMAX1DataOut_F1_106  ,
 REGofMAX1DataOut_F1_122, REGofMAX1DataOut_F1_124 , REGofMAX1DataOut_F1_126 , REGofMAX1DataOut_F1_128 , REGofMAX1DataOut_F1_130 , bigaddress222, Super_3_2_1_2_ch1 );
SUPERMUXMODULECONV2_new mux3_3_1_2_ch1 ( REGofMAX1DataOut_F1_27, REGofMAX1DataOut_F1_29 , REGofMAX1DataOut_F1_31 , REGofMAX1DataOut_F1_33 , REGofMAX1DataOut_F1_35 , REGofMAX1DataOut_F1_51 ,
REGofMAX1DataOut_F1_53 , REGofMAX1DataOut_F1_55 , REGofMAX1DataOut_F1_57 , REGofMAX1DataOut_F1_59 , REGofMAX1DataOut_F1_75 , REGofMAX1DataOut_F1_77 , REGofMAX1DataOut_F1_79 ,
 REGofMAX1DataOut_F1_81 , REGofMAX1DataOut_F1_83 ,REGofMAX1DataOut_F1_99  , REGofMAX1DataOut_F1_101 , REGofMAX1DataOut_F1_103 , REGofMAX1DataOut_F1_105 , REGofMAX1DataOut_F1_107 ,
 REGofMAX1DataOut_F1_123, REGofMAX1DataOut_F1_125 , REGofMAX1DataOut_F1_127 , REGofMAX1DataOut_F1_129 , REGofMAX1DataOut_F1_131 , bigaddress222, Super_3_3_1_2_ch1 );


SUPERMUXMODULECONV2_new mux1_1_2_1_ch1 ( REGofMAX1DataOut_F1_12, REGofMAX1DataOut_F1_14 , REGofMAX1DataOut_F1_16 , REGofMAX1DataOut_F1_18 , REGofMAX1DataOut_F1_20 , REGofMAX1DataOut_F1_36 ,
 REGofMAX1DataOut_F1_38 , REGofMAX1DataOut_F1_40 , REGofMAX1DataOut_F1_42 , REGofMAX1DataOut_F1_44 , REGofMAX1DataOut_F1_60 , REGofMAX1DataOut_F1_62 , REGofMAX1DataOut_F1_64 ,
 REGofMAX1DataOut_F1_66, REGofMAX1DataOut_F1_68 , REGofMAX1DataOut_F1_84 , REGofMAX1DataOut_F1_86 , REGofMAX1DataOut_F1_88 , REGofMAX1DataOut_F1_90 , REGofMAX1DataOut_F1_92 ,
 REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_110  , REGofMAX1DataOut_F1_112 , REGofMAX1DataOut_F1_114 , REGofMAX1DataOut_F1_116 , bigaddress222, Super_1_1_2_1_ch1 );
SUPERMUXMODULECONV2_new mux1_2_2_1_ch1 ( REGofMAX1DataOut_F1_13, REGofMAX1DataOut_F1_15 , REGofMAX1DataOut_F1_17 , REGofMAX1DataOut_F1_19 , REGofMAX1DataOut_F1_21 , REGofMAX1DataOut_F1_37 ,
 REGofMAX1DataOut_F1_39 , REGofMAX1DataOut_F1_41 , REGofMAX1DataOut_F1_43 , REGofMAX1DataOut_F1_45 , REGofMAX1DataOut_F1_61 , REGofMAX1DataOut_F1_63 , REGofMAX1DataOut_F1_65 ,
 REGofMAX1DataOut_F1_67, REGofMAX1DataOut_F1_69 , REGofMAX1DataOut_F1_85 , REGofMAX1DataOut_F1_87 , REGofMAX1DataOut_F1_89 , REGofMAX1DataOut_F1_91 , REGofMAX1DataOut_F1_93 ,
 REGofMAX1DataOut_F1_109, REGofMAX1DataOut_F1_111 , REGofMAX1DataOut_F1_113 , REGofMAX1DataOut_F1_115 , REGofMAX1DataOut_F1_117 , bigaddress222, Super_1_2_2_1_ch1 );
SUPERMUXMODULECONV2_new mux1_3_2_1_ch1 ( REGofMAX1DataOut_F1_14, REGofMAX1DataOut_F1_16 , REGofMAX1DataOut_F1_18 , REGofMAX1DataOut_F1_20 , REGofMAX1DataOut_F1_22 , REGofMAX1DataOut_F1_38 ,
REGofMAX1DataOut_F1_40  , REGofMAX1DataOut_F1_42 , REGofMAX1DataOut_F1_44 , REGofMAX1DataOut_F1_46 , REGofMAX1DataOut_F1_62 , REGofMAX1DataOut_F1_64 ,REGofMAX1DataOut_F1_66 ,
 REGofMAX1DataOut_F1_68 , REGofMAX1DataOut_F1_70 , REGofMAX1DataOut_F1_86 , REGofMAX1DataOut_F1_88 ,REGofMAX1DataOut_F1_90  , REGofMAX1DataOut_F1_92 , REGofMAX1DataOut_F1_94 ,
REGofMAX1DataOut_F1_110 , REGofMAX1DataOut_F1_112 , REGofMAX1DataOut_F1_114 , REGofMAX1DataOut_F1_116 , REGofMAX1DataOut_F1_118 , bigaddress222, Super_1_3_2_1_ch1 );
SUPERMUXMODULECONV2_new mux2_1_2_1_ch1 ( REGofMAX1DataOut_F1_24, REGofMAX1DataOut_F1_26 , REGofMAX1DataOut_F1_28 , REGofMAX1DataOut_F1_30 , REGofMAX1DataOut_F1_32 , REGofMAX1DataOut_F1_48 ,
 REGofMAX1DataOut_F1_50 , REGofMAX1DataOut_F1_52 , REGofMAX1DataOut_F1_54 , REGofMAX1DataOut_F1_56 , REGofMAX1DataOut_F1_72 , REGofMAX1DataOut_F1_74 ,REGofMAX1DataOut_F1_76  ,
 REGofMAX1DataOut_F1_78, REGofMAX1DataOut_F1_80 , REGofMAX1DataOut_F1_96 , REGofMAX1DataOut_F1_98 , REGofMAX1DataOut_F1_100 , REGofMAX1DataOut_F1_102 , REGofMAX1DataOut_F1_104 ,
REGofMAX1DataOut_F1_120 , REGofMAX1DataOut_F1_122 , REGofMAX1DataOut_F1_124 , REGofMAX1DataOut_F1_126 , REGofMAX1DataOut_F1_128 , bigaddress222, Super_2_1_2_1_ch1 );
SUPERMUXMODULECONV2_new mux2_2_2_1_ch1 ( REGofMAX1DataOut_F1_25, REGofMAX1DataOut_F1_27 , REGofMAX1DataOut_F1_29 , REGofMAX1DataOut_F1_31 , REGofMAX1DataOut_F1_33 , REGofMAX1DataOut_F1_49 ,
 REGofMAX1DataOut_F1_51 , REGofMAX1DataOut_F1_53 , REGofMAX1DataOut_F1_55 , REGofMAX1DataOut_F1_57 , REGofMAX1DataOut_F1_73 , REGofMAX1DataOut_F1_75 , REGofMAX1DataOut_F1_77 ,
 REGofMAX1DataOut_F1_79, REGofMAX1DataOut_F1_81 , REGofMAX1DataOut_F1_97 , REGofMAX1DataOut_F1_99 , REGofMAX1DataOut_F1_101 , REGofMAX1DataOut_F1_103 , REGofMAX1DataOut_F1_105 ,
REGofMAX1DataOut_F1_121 , REGofMAX1DataOut_F1_123 , REGofMAX1DataOut_F1_125 , REGofMAX1DataOut_F1_127 , REGofMAX1DataOut_F1_129 , bigaddress222, Super_2_2_2_1_ch1 );
SUPERMUXMODULECONV2_new mux2_3_2_1_ch1 ( REGofMAX1DataOut_F1_26, REGofMAX1DataOut_F1_28 , REGofMAX1DataOut_F1_30 , REGofMAX1DataOut_F1_32 , REGofMAX1DataOut_F1_34 , REGofMAX1DataOut_F1_50 ,
 REGofMAX1DataOut_F1_52 , REGofMAX1DataOut_F1_54 , REGofMAX1DataOut_F1_56 , REGofMAX1DataOut_F1_58 , REGofMAX1DataOut_F1_74 , REGofMAX1DataOut_F1_76 ,REGofMAX1DataOut_F1_78  ,
 REGofMAX1DataOut_F1_80, REGofMAX1DataOut_F1_82 , REGofMAX1DataOut_F1_98 , REGofMAX1DataOut_F1_100 , REGofMAX1DataOut_F1_102 , REGofMAX1DataOut_F1_104 , REGofMAX1DataOut_F1_106 ,
 REGofMAX1DataOut_F1_122, REGofMAX1DataOut_F1_124 , REGofMAX1DataOut_F1_126 , REGofMAX1DataOut_F1_128 , REGofMAX1DataOut_F1_130 , bigaddress222, Super_2_3_2_1_ch1 );
SUPERMUXMODULECONV2_new mux3_1_2_1_ch1 ( REGofMAX1DataOut_F1_36, REGofMAX1DataOut_F1_38 , REGofMAX1DataOut_F1_40 , REGofMAX1DataOut_F1_42 , REGofMAX1DataOut_F1_44 , REGofMAX1DataOut_F1_60 ,
 REGofMAX1DataOut_F1_62 , REGofMAX1DataOut_F1_64 , REGofMAX1DataOut_F1_66 , REGofMAX1DataOut_F1_68 , REGofMAX1DataOut_F1_84 , REGofMAX1DataOut_F1_86 ,REGofMAX1DataOut_F1_88  ,
 REGofMAX1DataOut_F1_90, REGofMAX1DataOut_F1_92 , REGofMAX1DataOut_F1_108 , REGofMAX1DataOut_F1_110 , REGofMAX1DataOut_F1_112 , REGofMAX1DataOut_F1_114 , REGofMAX1DataOut_F1_116 ,
 REGofMAX1DataOut_F1_132, REGofMAX1DataOut_F1_134 , REGofMAX1DataOut_F1_136 , REGofMAX1DataOut_F1_138 , REGofMAX1DataOut_F1_140 , bigaddress222, Super_3_1_2_1_ch1 );
SUPERMUXMODULECONV2_new mux3_2_2_1_ch1 ( REGofMAX1DataOut_F1_37, REGofMAX1DataOut_F1_39 , REGofMAX1DataOut_F1_41 , REGofMAX1DataOut_F1_43 , REGofMAX1DataOut_F1_45 , REGofMAX1DataOut_F1_61 ,
 REGofMAX1DataOut_F1_63 , REGofMAX1DataOut_F1_65 , REGofMAX1DataOut_F1_67 , REGofMAX1DataOut_F1_69 , REGofMAX1DataOut_F1_85 , REGofMAX1DataOut_F1_87 , REGofMAX1DataOut_F1_89 ,
 REGofMAX1DataOut_F1_91, REGofMAX1DataOut_F1_93 , REGofMAX1DataOut_F1_109 , REGofMAX1DataOut_F1_111 , REGofMAX1DataOut_F1_113 , REGofMAX1DataOut_F1_115 , REGofMAX1DataOut_F1_117 ,
 REGofMAX1DataOut_F1_133, REGofMAX1DataOut_F1_135 , REGofMAX1DataOut_F1_137 , REGofMAX1DataOut_F1_139 , REGofMAX1DataOut_F1_141 , bigaddress222, Super_3_2_2_1_ch1 );
SUPERMUXMODULECONV2_new mux3_3_2_1_ch1 ( REGofMAX1DataOut_F1_38, REGofMAX1DataOut_F1_40 , REGofMAX1DataOut_F1_42 , REGofMAX1DataOut_F1_44 , REGofMAX1DataOut_F1_46 , REGofMAX1DataOut_F1_62 ,
 REGofMAX1DataOut_F1_64 , REGofMAX1DataOut_F1_66 , REGofMAX1DataOut_F1_68 , REGofMAX1DataOut_F1_70 , REGofMAX1DataOut_F1_86 , REGofMAX1DataOut_F1_88 , REGofMAX1DataOut_F1_90 ,
 REGofMAX1DataOut_F1_92, REGofMAX1DataOut_F1_94 , REGofMAX1DataOut_F1_110 , REGofMAX1DataOut_F1_112 , REGofMAX1DataOut_F1_114 , REGofMAX1DataOut_F1_116 , REGofMAX1DataOut_F1_118 ,
 REGofMAX1DataOut_F1_134,  REGofMAX1DataOut_F1_136, REGofMAX1DataOut_F1_138 , REGofMAX1DataOut_F1_140 , REGofMAX1DataOut_F1_142 , bigaddress222, Super_3_3_2_1_ch1 );


SUPERMUXMODULECONV2_new mux1_1_2_2_ch1 ( REGofMAX1DataOut_F1_13, REGofMAX1DataOut_F1_15 , REGofMAX1DataOut_F1_17 , REGofMAX1DataOut_F1_19 , REGofMAX1DataOut_F1_21 , REGofMAX1DataOut_F1_37 ,
 REGofMAX1DataOut_F1_39 , REGofMAX1DataOut_F1_41 , REGofMAX1DataOut_F1_43 , REGofMAX1DataOut_F1_45 , REGofMAX1DataOut_F1_61 , REGofMAX1DataOut_F1_63 , REGofMAX1DataOut_F1_65 ,
 REGofMAX1DataOut_F1_67, REGofMAX1DataOut_F1_69 , REGofMAX1DataOut_F1_85 , REGofMAX1DataOut_F1_87 , REGofMAX1DataOut_F1_89 , REGofMAX1DataOut_F1_91 , REGofMAX1DataOut_F1_93 ,
 REGofMAX1DataOut_F1_109, REGofMAX1DataOut_F1_111 , REGofMAX1DataOut_F1_113 , REGofMAX1DataOut_F1_115 , REGofMAX1DataOut_F1_117 , bigaddress222, Super_1_1_2_2_ch1 );
SUPERMUXMODULECONV2_new mux1_2_2_2_ch1 ( REGofMAX1DataOut_F1_14, REGofMAX1DataOut_F1_16 , REGofMAX1DataOut_F1_18 , REGofMAX1DataOut_F1_20 , REGofMAX1DataOut_F1_22 , REGofMAX1DataOut_F1_38 ,
 REGofMAX1DataOut_F1_40 , REGofMAX1DataOut_F1_42 , REGofMAX1DataOut_F1_44 , REGofMAX1DataOut_F1_46 , REGofMAX1DataOut_F1_62 , REGofMAX1DataOut_F1_64 , REGofMAX1DataOut_F1_66 ,
REGofMAX1DataOut_F1_68 , REGofMAX1DataOut_F1_70 , REGofMAX1DataOut_F1_86 , REGofMAX1DataOut_F1_88 , REGofMAX1DataOut_F1_90 , REGofMAX1DataOut_F1_92 , REGofMAX1DataOut_F1_94 ,
 REGofMAX1DataOut_F1_110 , REGofMAX1DataOut_F1_112 , REGofMAX1DataOut_F1_114 , REGofMAX1DataOut_F1_116 , REGofMAX1DataOut_F1_118 , bigaddress222, Super_1_2_2_2_ch1 );
SUPERMUXMODULECONV2_new mux1_3_2_2_ch1 ( REGofMAX1DataOut_F1_15, REGofMAX1DataOut_F1_17 , REGofMAX1DataOut_F1_19 , REGofMAX1DataOut_F1_21 , REGofMAX1DataOut_F1_23 , REGofMAX1DataOut_F1_39 ,
 REGofMAX1DataOut_F1_41 , REGofMAX1DataOut_F1_43 , REGofMAX1DataOut_F1_45 , REGofMAX1DataOut_F1_47 , REGofMAX1DataOut_F1_63 , REGofMAX1DataOut_F1_65 , REGofMAX1DataOut_F1_67 ,
 REGofMAX1DataOut_F1_69, REGofMAX1DataOut_F1_71 , REGofMAX1DataOut_F1_87 , REGofMAX1DataOut_F1_89 , REGofMAX1DataOut_F1_91 , REGofMAX1DataOut_F1_93 , REGofMAX1DataOut_F1_95 ,
 REGofMAX1DataOut_F1_111, REGofMAX1DataOut_F1_113 , REGofMAX1DataOut_F1_115 , REGofMAX1DataOut_F1_117 , REGofMAX1DataOut_F1_119 , bigaddress222, Super_1_3_2_2_ch1 );
SUPERMUXMODULECONV2_new mux2_1_2_2_ch1 ( REGofMAX1DataOut_F1_25, REGofMAX1DataOut_F1_27 , REGofMAX1DataOut_F1_29 , REGofMAX1DataOut_F1_31 , REGofMAX1DataOut_F1_33 , REGofMAX1DataOut_F1_49 ,
 REGofMAX1DataOut_F1_51 , REGofMAX1DataOut_F1_53 , REGofMAX1DataOut_F1_55 , REGofMAX1DataOut_F1_57 , REGofMAX1DataOut_F1_73 , REGofMAX1DataOut_F1_75 , REGofMAX1DataOut_F1_77 ,
 REGofMAX1DataOut_F1_79, REGofMAX1DataOut_F1_81 , REGofMAX1DataOut_F1_97 , REGofMAX1DataOut_F1_99 , REGofMAX1DataOut_F1_101 , REGofMAX1DataOut_F1_103 , REGofMAX1DataOut_F1_105 ,
 REGofMAX1DataOut_F1_121, REGofMAX1DataOut_F1_123 , REGofMAX1DataOut_F1_125 , REGofMAX1DataOut_F1_127 , REGofMAX1DataOut_F1_129 , bigaddress222, Super_2_1_2_2_ch1 );
SUPERMUXMODULECONV2_new mux2_2_2_2_ch1 ( REGofMAX1DataOut_F1_26, REGofMAX1DataOut_F1_28 , REGofMAX1DataOut_F1_30 , REGofMAX1DataOut_F1_32 , REGofMAX1DataOut_F1_34 , REGofMAX1DataOut_F1_50 ,
 REGofMAX1DataOut_F1_52 , REGofMAX1DataOut_F1_54 , REGofMAX1DataOut_F1_56 , REGofMAX1DataOut_F1_58 , REGofMAX1DataOut_F1_74 , REGofMAX1DataOut_F1_76 , REGofMAX1DataOut_F1_78 ,
 REGofMAX1DataOut_F1_80, REGofMAX1DataOut_F1_82 , REGofMAX1DataOut_F1_98 , REGofMAX1DataOut_F1_100 , REGofMAX1DataOut_F1_102 , REGofMAX1DataOut_F1_104 , REGofMAX1DataOut_F1_106 ,
 REGofMAX1DataOut_F1_122, REGofMAX1DataOut_F1_124 , REGofMAX1DataOut_F1_126 , REGofMAX1DataOut_F1_128 , REGofMAX1DataOut_F1_130 , bigaddress222, Super_2_2_2_2_ch1 );
SUPERMUXMODULECONV2_new mux2_3_2_2_ch1 ( REGofMAX1DataOut_F1_27, REGofMAX1DataOut_F1_29 , REGofMAX1DataOut_F1_31 , REGofMAX1DataOut_F1_33 , REGofMAX1DataOut_F1_35 , REGofMAX1DataOut_F1_51 ,
 REGofMAX1DataOut_F1_53 , REGofMAX1DataOut_F1_55 , REGofMAX1DataOut_F1_57 , REGofMAX1DataOut_F1_59 , REGofMAX1DataOut_F1_75 , REGofMAX1DataOut_F1_77 , REGofMAX1DataOut_F1_79 ,
 REGofMAX1DataOut_F1_81, REGofMAX1DataOut_F1_83 , REGofMAX1DataOut_F1_99 , REGofMAX1DataOut_F1_101 , REGofMAX1DataOut_F1_103 , REGofMAX1DataOut_F1_105 , REGofMAX1DataOut_F1_107 ,
 REGofMAX1DataOut_F1_123, REGofMAX1DataOut_F1_125 , REGofMAX1DataOut_F1_127 , REGofMAX1DataOut_F1_129 , REGofMAX1DataOut_F1_131 , bigaddress222, Super_2_3_2_2_ch1 );
SUPERMUXMODULECONV2_new mux3_1_2_2_ch1 ( REGofMAX1DataOut_F1_37, REGofMAX1DataOut_F1_39 , REGofMAX1DataOut_F1_41 , REGofMAX1DataOut_F1_43 , REGofMAX1DataOut_F1_45 , REGofMAX1DataOut_F1_61 ,
 REGofMAX1DataOut_F1_63 , REGofMAX1DataOut_F1_65 , REGofMAX1DataOut_F1_67 , REGofMAX1DataOut_F1_69 , REGofMAX1DataOut_F1_85 , REGofMAX1DataOut_F1_87 , REGofMAX1DataOut_F1_89 ,
 REGofMAX1DataOut_F1_91, REGofMAX1DataOut_F1_93 , REGofMAX1DataOut_F1_109 , REGofMAX1DataOut_F1_111 , REGofMAX1DataOut_F1_113 , REGofMAX1DataOut_F1_115 , REGofMAX1DataOut_F1_117 ,
 REGofMAX1DataOut_F1_133, REGofMAX1DataOut_F1_135 ,REGofMAX1DataOut_F1_137  , REGofMAX1DataOut_F1_139 , REGofMAX1DataOut_F1_141 , bigaddress222, Super_3_1_2_2_ch1 );
SUPERMUXMODULECONV2_new mux3_2_2_2_ch1 ( REGofMAX1DataOut_F1_38, REGofMAX1DataOut_F1_40 , REGofMAX1DataOut_F1_42 , REGofMAX1DataOut_F1_44 , REGofMAX1DataOut_F1_46 , REGofMAX1DataOut_F1_62 ,
 REGofMAX1DataOut_F1_64 , REGofMAX1DataOut_F1_66 , REGofMAX1DataOut_F1_68 , REGofMAX1DataOut_F1_70 , REGofMAX1DataOut_F1_86 , REGofMAX1DataOut_F1_88 , REGofMAX1DataOut_F1_90 ,
 REGofMAX1DataOut_F1_92, REGofMAX1DataOut_F1_94 , REGofMAX1DataOut_F1_110 , REGofMAX1DataOut_F1_112 , REGofMAX1DataOut_F1_114 , REGofMAX1DataOut_F1_116 , REGofMAX1DataOut_F1_118 ,
REGofMAX1DataOut_F1_134 , REGofMAX1DataOut_F1_136 , REGofMAX1DataOut_F1_138 , REGofMAX1DataOut_F1_140 , REGofMAX1DataOut_F1_142 , bigaddress222, Super_3_2_2_2_ch1 );
SUPERMUXMODULECONV2_new mux3_3_2_2_ch1 ( REGofMAX1DataOut_F1_39, REGofMAX1DataOut_F1_41 , REGofMAX1DataOut_F1_43 , REGofMAX1DataOut_F1_45 , REGofMAX1DataOut_F1_47 , REGofMAX1DataOut_F1_63 ,
 REGofMAX1DataOut_F1_65 , REGofMAX1DataOut_F1_67 , REGofMAX1DataOut_F1_69 , REGofMAX1DataOut_F1_71 , REGofMAX1DataOut_F1_87 , REGofMAX1DataOut_F1_89 , REGofMAX1DataOut_F1_91 ,
 REGofMAX1DataOut_F1_93, REGofMAX1DataOut_F1_95 , REGofMAX1DataOut_F1_111 , REGofMAX1DataOut_F1_113 , REGofMAX1DataOut_F1_115 , REGofMAX1DataOut_F1_117 , REGofMAX1DataOut_F1_119 ,
 REGofMAX1DataOut_F1_135, REGofMAX1DataOut_F1_137 , REGofMAX1DataOut_F1_139 , REGofMAX1DataOut_F1_141 ,  REGofMAX1DataOut_F1_143, bigaddress222, Super_3_3_2_2_ch1 );


MUX9X1_conv2 CONV2_MUX0 ( Super_1_1_1_1_ch1 , Super_1_2_1_1_ch1 , Super_1_3_1_1_ch1 , Super_2_1_1_1_ch1 , Super_2_2_1_1_ch1 , Super_2_3_1_1_ch1 , Super_3_1_1_1_ch1 , Super_3_2_1_1_ch1 , Super_3_3_1_1_ch1 ,  CONV2_address , In1_CONV2_MUXout0 );
MUX9X1_conv2 CONV2_MUX1 ( Super_1_1_1_2_ch1 , Super_1_2_1_2_ch1 , Super_1_3_1_2_ch1 , Super_2_1_1_2_ch1 , Super_2_2_1_2_ch1 , Super_2_3_1_2_ch1 , Super_3_1_1_2_ch1 , Super_3_2_1_2_ch1 , Super_3_3_1_2_ch1 ,  CONV2_address , In1_CONV2_MUXout1 );
MUX9X1_conv2 CONV2_MUX10 ( Super_1_1_2_1_ch1 , Super_1_2_2_1_ch1 , Super_1_3_2_1_ch1 , Super_2_1_2_1_ch1 , Super_2_2_2_1_ch1 , Super_2_3_2_1_ch1 , Super_3_1_2_1_ch1 , Super_3_2_2_1_ch1 , Super_3_3_2_1_ch1 ,  CONV2_address , In1_CONV2_MUXout10 );
MUX9X1_conv2 CONV2_MUX11 ( Super_1_1_2_2_ch1 , Super_1_2_2_2_ch1 , Super_1_3_2_2_ch1 , Super_2_1_2_2_ch1 , Super_2_2_2_2_ch1 , Super_2_3_2_2_ch1 , Super_3_1_2_2_ch1 , Super_3_2_2_2_ch1 , Super_3_3_2_2_ch1 ,  CONV2_address , In1_CONV2_MUXout11 );



MAC_9 In1_CONV2_MAC0_F1 (In1_CONV2_ROMout, In1_CONV2_MUXout0 , clk, In1_CONV2_MACoutF1_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC1_F1  (In1_CONV2_ROMout, In1_CONV2_MUXout1 , clk, In1_CONV2_MACoutF1_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC10_F1  (In1_CONV2_ROMout, In1_CONV2_MUXout10 , clk, In1_CONV2_MACoutF1_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC11_F1  (In1_CONV2_ROMout, In1_CONV2_MUXout11 , clk, In1_CONV2_MACoutF1_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In1_CONV2_MAC0_F2 (In1_CONV2_ROMout1, In1_CONV2_MUXout0 , clk, In1_CONV2_MACoutF2_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC1_F2  (In1_CONV2_ROMout1, In1_CONV2_MUXout1 , clk, In1_CONV2_MACoutF2_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC10_F2  (In1_CONV2_ROMout1, In1_CONV2_MUXout10 , clk, In1_CONV2_MACoutF2_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC11_F2  (In1_CONV2_ROMout1, In1_CONV2_MUXout11 , clk, In1_CONV2_MACoutF2_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In1_CONV2_MAC0_F3 (In1_CONV2_ROMout2, In1_CONV2_MUXout0 , clk, In1_CONV2_MACoutF3_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC1_F3 (In1_CONV2_ROMout2, In1_CONV2_MUXout1 , clk, In1_CONV2_MACoutF3_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC10_F3 (In1_CONV2_ROMout2, In1_CONV2_MUXout10 , clk, In1_CONV2_MACoutF3_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC11_F3 (In1_CONV2_ROMout2, In1_CONV2_MUXout11 , clk, In1_CONV2_MACoutF3_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In1_CONV2_MAC0_F4 (In1_CONV2_ROMout3, In1_CONV2_MUXout0 , clk, In1_CONV2_MACoutF4_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC1_F4  (In1_CONV2_ROMout3, In1_CONV2_MUXout1 , clk, In1_CONV2_MACoutF4_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC10_F4  (In1_CONV2_ROMout3, In1_CONV2_MUXout10 , clk, In1_CONV2_MACoutF4_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In1_CONV2_MAC11_F4  (In1_CONV2_ROMout3, In1_CONV2_MUXout11 , clk, In1_CONV2_MACoutF4_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);



///2nd input channel

SUPERMUXMODULECONV2_new mux1_1_1_1_ch2 ( REGofMAX1DataOut_F2_0, REGofMAX1DataOut_F2_2 , REGofMAX1DataOut_F2_4 , REGofMAX1DataOut_F2_6 , REGofMAX1DataOut_F2_8 , REGofMAX1DataOut_F2_24 ,
 REGofMAX1DataOut_F2_26 , REGofMAX1DataOut_F2_28 , REGofMAX1DataOut_F2_30 , REGofMAX1DataOut_F2_32 , REGofMAX1DataOut_F2_48 , REGofMAX1DataOut_F2_50 , REGofMAX1DataOut_F2_52 ,
 REGofMAX1DataOut_F2_54, REGofMAX1DataOut_F2_56 , REGofMAX1DataOut_F2_72 , REGofMAX1DataOut_F2_74 , REGofMAX1DataOut_F2_76 , REGofMAX1DataOut_F2_78 , REGofMAX1DataOut_F2_80 ,
 REGofMAX1DataOut_F2_96, REGofMAX1DataOut_F2_98 ,REGofMAX1DataOut_F2_100  , REGofMAX1DataOut_F2_102 , REGofMAX1DataOut_F2_104 , bigaddress222, Super_1_1_1_1_ch2 );
SUPERMUXMODULECONV2_new mux1_2_1_1_ch2 ( REGofMAX1DataOut_F2_1 , REGofMAX1DataOut_F2_3 , REGofMAX1DataOut_F2_5 , REGofMAX1DataOut_F2_7 , REGofMAX1DataOut_F2_9 , REGofMAX1DataOut_F2_25 ,
 REGofMAX1DataOut_F2_27 , REGofMAX1DataOut_F2_29 , REGofMAX1DataOut_F2_31 , REGofMAX1DataOut_F2_33 , REGofMAX1DataOut_F2_49 , REGofMAX1DataOut_F2_51 , REGofMAX1DataOut_F2_53 ,
 REGofMAX1DataOut_F2_55, REGofMAX1DataOut_F2_57 , REGofMAX1DataOut_F2_73 , REGofMAX1DataOut_F2_75 , REGofMAX1DataOut_F2_77 , REGofMAX1DataOut_F2_79 , REGofMAX1DataOut_F2_81 ,
 REGofMAX1DataOut_F2_97, REGofMAX1DataOut_F2_99 , REGofMAX1DataOut_F2_101 , REGofMAX1DataOut_F2_103 ,  REGofMAX1DataOut_F2_105, bigaddress222, Super_1_2_1_1_ch2 );
SUPERMUXMODULECONV2_new mux1_3_1_1_ch2 ( REGofMAX1DataOut_F2_2,  REGofMAX1DataOut_F2_4, REGofMAX1DataOut_F2_6 , REGofMAX1DataOut_F2_8 , REGofMAX1DataOut_F2_10 , REGofMAX1DataOut_F2_26 ,
 REGofMAX1DataOut_F2_28 , REGofMAX1DataOut_F2_30 , REGofMAX1DataOut_F2_32 , REGofMAX1DataOut_F2_34 , REGofMAX1DataOut_F2_50 , REGofMAX1DataOut_F2_52 , REGofMAX1DataOut_F2_54 ,
 REGofMAX1DataOut_F2_56, REGofMAX1DataOut_F2_58 , REGofMAX1DataOut_F2_74 , REGofMAX1DataOut_F2_76 , REGofMAX1DataOut_F2_78 , REGofMAX1DataOut_F2_80 , REGofMAX1DataOut_F2_82 ,
 REGofMAX1DataOut_F2_98, REGofMAX1DataOut_F2_100 , REGofMAX1DataOut_F2_102 , REGofMAX1DataOut_F2_104 , REGofMAX1DataOut_F2_106 , bigaddress222, Super_1_3_1_1_ch2 );
SUPERMUXMODULECONV2_new mux2_1_1_1_ch2 ( REGofMAX1DataOut_F2_12 ,REGofMAX1DataOut_F2_14  , REGofMAX1DataOut_F2_16 , REGofMAX1DataOut_F2_18 , REGofMAX1DataOut_F2_20 , REGofMAX1DataOut_F2_36 ,
 REGofMAX1DataOut_F2_38 , REGofMAX1DataOut_F2_40 , REGofMAX1DataOut_F2_42 , REGofMAX1DataOut_F2_44 , REGofMAX1DataOut_F2_60 , REGofMAX1DataOut_F2_62 , REGofMAX1DataOut_F2_64 ,
 REGofMAX1DataOut_F2_66, REGofMAX1DataOut_F2_68 , REGofMAX1DataOut_F2_84 , REGofMAX1DataOut_F2_86 , REGofMAX1DataOut_F2_88 , REGofMAX1DataOut_F2_90 , REGofMAX1DataOut_F2_92  ,
 REGofMAX1DataOut_F2_108, REGofMAX1DataOut_F2_110 , REGofMAX1DataOut_F2_112 , REGofMAX1DataOut_F2_114 , REGofMAX1DataOut_F2_116 , bigaddress222, Super_2_1_1_1_ch2 );
SUPERMUXMODULECONV2_new mux2_2_1_1_ch2 ( REGofMAX1DataOut_F2_13, REGofMAX1DataOut_F2_15 , REGofMAX1DataOut_F2_17 , REGofMAX1DataOut_F2_19 , REGofMAX1DataOut_F2_21 , REGofMAX1DataOut_F2_37 ,
 REGofMAX1DataOut_F2_39 , REGofMAX1DataOut_F2_41 , REGofMAX1DataOut_F2_43 , REGofMAX1DataOut_F2_45 , REGofMAX1DataOut_F2_61 , REGofMAX1DataOut_F2_63 , REGofMAX1DataOut_F2_65 ,
 REGofMAX1DataOut_F2_67, REGofMAX1DataOut_F2_69 , REGofMAX1DataOut_F2_85 , REGofMAX1DataOut_F2_87 , REGofMAX1DataOut_F2_89 , REGofMAX1DataOut_F2_91 ,REGofMAX1DataOut_F2_93  ,
 REGofMAX1DataOut_F2_109, REGofMAX1DataOut_F2_111 , REGofMAX1DataOut_F2_113 , REGofMAX1DataOut_F2_115 ,REGofMAX1DataOut_F2_117  , bigaddress222, Super_2_2_1_1_ch2 );
SUPERMUXMODULECONV2_new mux2_3_1_1_ch2 ( REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_16  , REGofMAX1DataOut_F2_18 , REGofMAX1DataOut_F2_20 , REGofMAX1DataOut_F2_22 , REGofMAX1DataOut_F2_38 ,
 REGofMAX1DataOut_F2_40 , REGofMAX1DataOut_F2_42 , REGofMAX1DataOut_F2_44 , REGofMAX1DataOut_F2_46 , REGofMAX1DataOut_F2_62 , REGofMAX1DataOut_F2_64 , REGofMAX1DataOut_F2_66 ,
 REGofMAX1DataOut_F2_68, REGofMAX1DataOut_F2_70 , REGofMAX1DataOut_F2_86 , REGofMAX1DataOut_F2_88 , REGofMAX1DataOut_F2_90 , REGofMAX1DataOut_F2_92 , REGofMAX1DataOut_F2_94 ,
 REGofMAX1DataOut_F2_110, REGofMAX1DataOut_F2_112 , REGofMAX1DataOut_F2_114 , REGofMAX1DataOut_F2_116 , REGofMAX1DataOut_F2_118 , bigaddress222, Super_2_3_1_1_ch2 );
SUPERMUXMODULECONV2_new mux3_1_1_1_ch2 ( REGofMAX1DataOut_F2_24, REGofMAX1DataOut_F2_26 , REGofMAX1DataOut_F2_28 , REGofMAX1DataOut_F2_30 , REGofMAX1DataOut_F2_32 , REGofMAX1DataOut_F2_48 ,
 REGofMAX1DataOut_F2_50 , REGofMAX1DataOut_F2_52 , REGofMAX1DataOut_F2_54 , REGofMAX1DataOut_F2_56 , REGofMAX1DataOut_F2_72 , REGofMAX1DataOut_F2_74 , REGofMAX1DataOut_F2_76 ,
 REGofMAX1DataOut_F2_78, REGofMAX1DataOut_F2_80 , REGofMAX1DataOut_F2_96 , REGofMAX1DataOut_F2_98 , REGofMAX1DataOut_F2_100 , REGofMAX1DataOut_F2_102 , REGofMAX1DataOut_F2_104 ,
 REGofMAX1DataOut_F2_120, REGofMAX1DataOut_F2_122 , REGofMAX1DataOut_F2_124 , REGofMAX1DataOut_F2_126 , REGofMAX1DataOut_F2_128 , bigaddress222, Super_3_1_1_1_ch2 );
SUPERMUXMODULECONV2_new mux3_2_1_1_ch2 ( REGofMAX1DataOut_F2_25, REGofMAX1DataOut_F2_27 , REGofMAX1DataOut_F2_29 , REGofMAX1DataOut_F2_31 , REGofMAX1DataOut_F2_33 , REGofMAX1DataOut_F2_49 ,
 REGofMAX1DataOut_F2_51 ,REGofMAX1DataOut_F2_53  , REGofMAX1DataOut_F2_55 , REGofMAX1DataOut_F2_57 , REGofMAX1DataOut_F2_73 , REGofMAX1DataOut_F2_75 , REGofMAX1DataOut_F2_77 ,
REGofMAX1DataOut_F2_79 , REGofMAX1DataOut_F2_81 , REGofMAX1DataOut_F2_97 , REGofMAX1DataOut_F2_99 , REGofMAX1DataOut_F2_101 , REGofMAX1DataOut_F2_103 , REGofMAX1DataOut_F2_105 ,
 REGofMAX1DataOut_F2_121 , REGofMAX1DataOut_F2_123 , REGofMAX1DataOut_F2_125 , REGofMAX1DataOut_F2_127 , REGofMAX1DataOut_F2_129 , bigaddress222, Super_3_2_1_1_ch2 );
SUPERMUXMODULECONV2_new mux3_3_1_1_ch2 ( REGofMAX1DataOut_F2_26, REGofMAX1DataOut_F2_28 , REGofMAX1DataOut_F2_30 , REGofMAX1DataOut_F2_32 , REGofMAX1DataOut_F2_34 , REGofMAX1DataOut_F2_50 ,
REGofMAX1DataOut_F2_52  , REGofMAX1DataOut_F2_54 , REGofMAX1DataOut_F2_56 , REGofMAX1DataOut_F2_58 , REGofMAX1DataOut_F2_74 , REGofMAX1DataOut_F2_76 , REGofMAX1DataOut_F2_78 ,
REGofMAX1DataOut_F2_80 , REGofMAX1DataOut_F2_82 , REGofMAX1DataOut_F2_98 , REGofMAX1DataOut_F2_100 , REGofMAX1DataOut_F2_102 , REGofMAX1DataOut_F2_104 , REGofMAX1DataOut_F2_106 ,
 REGofMAX1DataOut_F2_122 , REGofMAX1DataOut_F2_124 , REGofMAX1DataOut_F2_126 , REGofMAX1DataOut_F2_128 , REGofMAX1DataOut_F2_130 , bigaddress222, Super_3_3_1_1_ch2 );



SUPERMUXMODULECONV2_new mux1_1_1_2_ch2 ( REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_3  , REGofMAX1DataOut_F2_5 , REGofMAX1DataOut_F2_7 , REGofMAX1DataOut_F2_9 , REGofMAX1DataOut_F2_25 ,
REGofMAX1DataOut_F2_27 , REGofMAX1DataOut_F2_29 , REGofMAX1DataOut_F2_31 , REGofMAX1DataOut_F2_33 , REGofMAX1DataOut_F2_49 , REGofMAX1DataOut_F2_51 ,REGofMAX1DataOut_F2_53  ,
 REGofMAX1DataOut_F2_55 ,REGofMAX1DataOut_F2_57  , REGofMAX1DataOut_F2_73 , REGofMAX1DataOut_F2_75 , REGofMAX1DataOut_F2_77 , REGofMAX1DataOut_F2_79 , REGofMAX1DataOut_F2_81 ,
 REGofMAX1DataOut_F2_97, REGofMAX1DataOut_F2_99 , REGofMAX1DataOut_F2_101 , REGofMAX1DataOut_F2_103 , REGofMAX1DataOut_F2_105 , bigaddress222, Super_1_1_1_2_ch2 );
SUPERMUXMODULECONV2_new mux1_2_1_2_ch2 ( REGofMAX1DataOut_F2_2, REGofMAX1DataOut_F2_4 , REGofMAX1DataOut_F2_6 , REGofMAX1DataOut_F2_8 , REGofMAX1DataOut_F2_10 , REGofMAX1DataOut_F2_26 ,
REGofMAX1DataOut_F2_28 , REGofMAX1DataOut_F2_30 , REGofMAX1DataOut_F2_32 , REGofMAX1DataOut_F2_34 , REGofMAX1DataOut_F2_50 , REGofMAX1DataOut_F2_52 ,REGofMAX1DataOut_F2_54  ,
 REGofMAX1DataOut_F2_56 , REGofMAX1DataOut_F2_58 , REGofMAX1DataOut_F2_74 , REGofMAX1DataOut_F2_76 , REGofMAX1DataOut_F2_78 , REGofMAX1DataOut_F2_80 , REGofMAX1DataOut_F2_82 ,
 REGofMAX1DataOut_F2_98, REGofMAX1DataOut_F2_100 , REGofMAX1DataOut_F2_102 , REGofMAX1DataOut_F2_104 , REGofMAX1DataOut_F2_106 , bigaddress222, Super_1_2_1_2_ch2 );
SUPERMUXMODULECONV2_new mux1_3_1_2_ch2 ( REGofMAX1DataOut_F2_3, REGofMAX1DataOut_F2_5 , REGofMAX1DataOut_F2_7 , REGofMAX1DataOut_F2_9 , REGofMAX1DataOut_F2_11 , REGofMAX1DataOut_F2_27 ,
REGofMAX1DataOut_F2_29 , REGofMAX1DataOut_F2_31 , REGofMAX1DataOut_F2_33 , REGofMAX1DataOut_F2_35 , REGofMAX1DataOut_F2_51 , REGofMAX1DataOut_F2_53 , REGofMAX1DataOut_F2_55 ,
 REGofMAX1DataOut_F2_57 , REGofMAX1DataOut_F2_59 , REGofMAX1DataOut_F2_75 , REGofMAX1DataOut_F2_77 , REGofMAX1DataOut_F2_79 , REGofMAX1DataOut_F2_81 , REGofMAX1DataOut_F2_83 ,
 REGofMAX1DataOut_F2_99, REGofMAX1DataOut_F2_101 , REGofMAX1DataOut_F2_103 , REGofMAX1DataOut_F2_105 , REGofMAX1DataOut_F2_107 , bigaddress222, Super_1_3_1_2_ch2 );
SUPERMUXMODULECONV2_new mux2_1_1_2_ch2 ( REGofMAX1DataOut_F2_13, REGofMAX1DataOut_F2_15 , REGofMAX1DataOut_F2_17 , REGofMAX1DataOut_F2_19 , REGofMAX1DataOut_F2_21 , REGofMAX1DataOut_F2_37 ,
REGofMAX1DataOut_F2_39 , REGofMAX1DataOut_F2_41 , REGofMAX1DataOut_F2_43 , REGofMAX1DataOut_F2_45 , REGofMAX1DataOut_F2_61 , REGofMAX1DataOut_F2_63  ,REGofMAX1DataOut_F2_65  ,
 REGofMAX1DataOut_F2_67 , REGofMAX1DataOut_F2_69 , REGofMAX1DataOut_F2_85 , REGofMAX1DataOut_F2_87 , REGofMAX1DataOut_F2_89 , REGofMAX1DataOut_F2_91 , REGofMAX1DataOut_F2_93 ,
 REGofMAX1DataOut_F2_109, REGofMAX1DataOut_F2_111 , REGofMAX1DataOut_F2_113 , REGofMAX1DataOut_F2_115 , REGofMAX1DataOut_F2_117 , bigaddress222, Super_2_1_1_2_ch2 );
SUPERMUXMODULECONV2_new mux2_2_1_2_ch2 ( REGofMAX1DataOut_F2_14, REGofMAX1DataOut_F2_16 , REGofMAX1DataOut_F2_18 , REGofMAX1DataOut_F2_20 , REGofMAX1DataOut_F2_22 , REGofMAX1DataOut_F2_38 ,
REGofMAX1DataOut_F2_40  , REGofMAX1DataOut_F2_42 , REGofMAX1DataOut_F2_44 , REGofMAX1DataOut_F2_46 , REGofMAX1DataOut_F2_62 , REGofMAX1DataOut_F2_64 ,REGofMAX1DataOut_F2_66  ,
 REGofMAX1DataOut_F2_68 , REGofMAX1DataOut_F2_70 , REGofMAX1DataOut_F2_86 , REGofMAX1DataOut_F2_88 , REGofMAX1DataOut_F2_90 , REGofMAX1DataOut_F2_92 , REGofMAX1DataOut_F2_94 ,
 REGofMAX1DataOut_F2_110, REGofMAX1DataOut_F2_112 , REGofMAX1DataOut_F2_114 , REGofMAX1DataOut_F2_116 , REGofMAX1DataOut_F2_118 , bigaddress222, Super_2_2_1_2_ch2 );
SUPERMUXMODULECONV2_new mux2_3_1_2_ch2 ( REGofMAX1DataOut_F2_15, REGofMAX1DataOut_F2_17 , REGofMAX1DataOut_F2_19 , REGofMAX1DataOut_F2_21 , REGofMAX1DataOut_F2_23 , REGofMAX1DataOut_F2_39 ,
REGofMAX1DataOut_F2_41  , REGofMAX1DataOut_F2_43 , REGofMAX1DataOut_F2_45 , REGofMAX1DataOut_F2_47 , REGofMAX1DataOut_F2_63 , REGofMAX1DataOut_F2_65 ,REGofMAX1DataOut_F2_67  ,
 REGofMAX1DataOut_F2_69 , REGofMAX1DataOut_F2_71 , REGofMAX1DataOut_F2_87 , REGofMAX1DataOut_F2_89 , REGofMAX1DataOut_F2_91 , REGofMAX1DataOut_F2_93 , REGofMAX1DataOut_F2_95 ,
 REGofMAX1DataOut_F2_111, REGofMAX1DataOut_F2_113 , REGofMAX1DataOut_F2_115 , REGofMAX1DataOut_F2_117 , REGofMAX1DataOut_F2_119 , bigaddress222, Super_2_3_1_2_ch2 );
SUPERMUXMODULECONV2_new mux3_1_1_2_ch2 ( REGofMAX1DataOut_F2_25, REGofMAX1DataOut_F2_27 , REGofMAX1DataOut_F2_29 , REGofMAX1DataOut_F2_31 , REGofMAX1DataOut_F2_33 , REGofMAX1DataOut_F2_49 ,
REGofMAX1DataOut_F2_51 , REGofMAX1DataOut_F2_53 , REGofMAX1DataOut_F2_55 , REGofMAX1DataOut_F2_57 , REGofMAX1DataOut_F2_73 , REGofMAX1DataOut_F2_75 ,REGofMAX1DataOut_F2_77  ,
 REGofMAX1DataOut_F2_79 , REGofMAX1DataOut_F2_81 , REGofMAX1DataOut_F2_97 , REGofMAX1DataOut_F2_99 , REGofMAX1DataOut_F2_101 , REGofMAX1DataOut_F2_103 , REGofMAX1DataOut_F2_105 ,
REGofMAX1DataOut_F2_121 , REGofMAX1DataOut_F2_123 , REGofMAX1DataOut_F2_125 , REGofMAX1DataOut_F2_127 , REGofMAX1DataOut_F2_129 , bigaddress222, Super_3_1_1_2_ch2 );
SUPERMUXMODULECONV2_new mux3_2_1_2_ch2 ( REGofMAX1DataOut_F2_26, REGofMAX1DataOut_F2_28 , REGofMAX1DataOut_F2_30 , REGofMAX1DataOut_F2_32 , REGofMAX1DataOut_F2_34 , REGofMAX1DataOut_F2_50 ,
REGofMAX1DataOut_F2_52  , REGofMAX1DataOut_F2_54 , REGofMAX1DataOut_F2_56 , REGofMAX1DataOut_F2_58 , REGofMAX1DataOut_F2_74 , REGofMAX1DataOut_F2_76 ,REGofMAX1DataOut_F2_78  ,
 REGofMAX1DataOut_F2_80 , REGofMAX1DataOut_F2_82 , REGofMAX1DataOut_F2_98 , REGofMAX1DataOut_F2_100 , REGofMAX1DataOut_F2_102 , REGofMAX1DataOut_F2_104 ,REGofMAX1DataOut_F2_106  ,
 REGofMAX1DataOut_F2_122, REGofMAX1DataOut_F2_124 , REGofMAX1DataOut_F2_126 , REGofMAX1DataOut_F2_128 , REGofMAX1DataOut_F2_130 , bigaddress222, Super_3_2_1_2_ch2 );
SUPERMUXMODULECONV2_new mux3_3_1_2_ch2 ( REGofMAX1DataOut_F2_27, REGofMAX1DataOut_F2_29 , REGofMAX1DataOut_F2_31 , REGofMAX1DataOut_F2_33 , REGofMAX1DataOut_F2_35 , REGofMAX1DataOut_F2_51 ,
REGofMAX1DataOut_F2_53 , REGofMAX1DataOut_F2_55 , REGofMAX1DataOut_F2_57 , REGofMAX1DataOut_F2_59 , REGofMAX1DataOut_F2_75 , REGofMAX1DataOut_F2_77 , REGofMAX1DataOut_F2_79 ,
 REGofMAX1DataOut_F2_81 , REGofMAX1DataOut_F2_83 ,REGofMAX1DataOut_F2_99  , REGofMAX1DataOut_F2_101 , REGofMAX1DataOut_F2_103 , REGofMAX1DataOut_F2_105 , REGofMAX1DataOut_F2_107 ,
 REGofMAX1DataOut_F2_123, REGofMAX1DataOut_F2_125 , REGofMAX1DataOut_F2_127 , REGofMAX1DataOut_F2_129 , REGofMAX1DataOut_F2_131 , bigaddress222, Super_3_3_1_2_ch2 );


SUPERMUXMODULECONV2_new mux1_1_2_1_ch2 ( REGofMAX1DataOut_F2_12, REGofMAX1DataOut_F2_14 , REGofMAX1DataOut_F2_16 , REGofMAX1DataOut_F2_18 , REGofMAX1DataOut_F2_20 , REGofMAX1DataOut_F2_36 ,
 REGofMAX1DataOut_F2_38 , REGofMAX1DataOut_F2_40 , REGofMAX1DataOut_F2_42 , REGofMAX1DataOut_F2_44 , REGofMAX1DataOut_F2_60 , REGofMAX1DataOut_F2_62 , REGofMAX1DataOut_F2_64 ,
 REGofMAX1DataOut_F2_66, REGofMAX1DataOut_F2_68 , REGofMAX1DataOut_F2_84 , REGofMAX1DataOut_F2_86 , REGofMAX1DataOut_F2_88 , REGofMAX1DataOut_F2_90 , REGofMAX1DataOut_F2_92 ,
 REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_110  , REGofMAX1DataOut_F2_112 , REGofMAX1DataOut_F2_114 , REGofMAX1DataOut_F2_116 , bigaddress222, Super_1_1_2_1_ch2 );
SUPERMUXMODULECONV2_new mux1_2_2_1_ch2 ( REGofMAX1DataOut_F2_13, REGofMAX1DataOut_F2_15 , REGofMAX1DataOut_F2_17 , REGofMAX1DataOut_F2_19 , REGofMAX1DataOut_F2_21 , REGofMAX1DataOut_F2_37 ,
 REGofMAX1DataOut_F2_39 , REGofMAX1DataOut_F2_41 , REGofMAX1DataOut_F2_43 , REGofMAX1DataOut_F2_45 , REGofMAX1DataOut_F2_61 , REGofMAX1DataOut_F2_63 , REGofMAX1DataOut_F2_65 ,
 REGofMAX1DataOut_F2_67, REGofMAX1DataOut_F2_69 , REGofMAX1DataOut_F2_85 , REGofMAX1DataOut_F2_87 , REGofMAX1DataOut_F2_89 , REGofMAX1DataOut_F2_91 , REGofMAX1DataOut_F2_93 ,
 REGofMAX1DataOut_F2_109, REGofMAX1DataOut_F2_111 , REGofMAX1DataOut_F2_113 , REGofMAX1DataOut_F2_115 , REGofMAX1DataOut_F2_117 , bigaddress222, Super_1_2_2_1_ch2 );
SUPERMUXMODULECONV2_new mux1_3_2_1_ch2 ( REGofMAX1DataOut_F2_14, REGofMAX1DataOut_F2_16 , REGofMAX1DataOut_F2_18 , REGofMAX1DataOut_F2_20 , REGofMAX1DataOut_F2_22 , REGofMAX1DataOut_F2_38 ,
REGofMAX1DataOut_F2_40  , REGofMAX1DataOut_F2_42 , REGofMAX1DataOut_F2_44 , REGofMAX1DataOut_F2_46 , REGofMAX1DataOut_F2_62 , REGofMAX1DataOut_F2_64 ,REGofMAX1DataOut_F2_66 ,
 REGofMAX1DataOut_F2_68 , REGofMAX1DataOut_F2_70 , REGofMAX1DataOut_F2_86 , REGofMAX1DataOut_F2_88 ,REGofMAX1DataOut_F2_90  , REGofMAX1DataOut_F2_92 , REGofMAX1DataOut_F2_94 ,
REGofMAX1DataOut_F2_110 , REGofMAX1DataOut_F2_112 , REGofMAX1DataOut_F2_114 , REGofMAX1DataOut_F2_116 , REGofMAX1DataOut_F2_118 , bigaddress222, Super_1_3_2_1_ch2 );
SUPERMUXMODULECONV2_new mux2_1_2_1_ch2 ( REGofMAX1DataOut_F2_24, REGofMAX1DataOut_F2_26 , REGofMAX1DataOut_F2_28 , REGofMAX1DataOut_F2_30 , REGofMAX1DataOut_F2_32 , REGofMAX1DataOut_F2_48 ,
 REGofMAX1DataOut_F2_50 , REGofMAX1DataOut_F2_52 , REGofMAX1DataOut_F2_54 , REGofMAX1DataOut_F2_56 , REGofMAX1DataOut_F2_72 , REGofMAX1DataOut_F2_74 ,REGofMAX1DataOut_F2_76  ,
 REGofMAX1DataOut_F2_78, REGofMAX1DataOut_F2_80 , REGofMAX1DataOut_F2_96 , REGofMAX1DataOut_F2_98 , REGofMAX1DataOut_F2_100 , REGofMAX1DataOut_F2_102 , REGofMAX1DataOut_F2_104 ,
REGofMAX1DataOut_F2_120 , REGofMAX1DataOut_F2_122 , REGofMAX1DataOut_F2_124 , REGofMAX1DataOut_F2_126 , REGofMAX1DataOut_F2_128 , bigaddress222, Super_2_1_2_1_ch2 );
SUPERMUXMODULECONV2_new mux2_2_2_1_ch2 ( REGofMAX1DataOut_F2_25, REGofMAX1DataOut_F2_27 , REGofMAX1DataOut_F2_29 , REGofMAX1DataOut_F2_31 , REGofMAX1DataOut_F2_33 , REGofMAX1DataOut_F2_49 ,
 REGofMAX1DataOut_F2_51 , REGofMAX1DataOut_F2_53 , REGofMAX1DataOut_F2_55 , REGofMAX1DataOut_F2_57 , REGofMAX1DataOut_F2_73 , REGofMAX1DataOut_F2_75 , REGofMAX1DataOut_F2_77 ,
 REGofMAX1DataOut_F2_79, REGofMAX1DataOut_F2_81 , REGofMAX1DataOut_F2_97 , REGofMAX1DataOut_F2_99 , REGofMAX1DataOut_F2_101 , REGofMAX1DataOut_F2_103 , REGofMAX1DataOut_F2_105 ,
REGofMAX1DataOut_F2_121 , REGofMAX1DataOut_F2_123 , REGofMAX1DataOut_F2_125 , REGofMAX1DataOut_F2_127 , REGofMAX1DataOut_F2_129 , bigaddress222, Super_2_2_2_1_ch2 );
SUPERMUXMODULECONV2_new mux2_3_2_1_ch2 ( REGofMAX1DataOut_F2_26, REGofMAX1DataOut_F2_28 , REGofMAX1DataOut_F2_30 , REGofMAX1DataOut_F2_32 , REGofMAX1DataOut_F2_34 , REGofMAX1DataOut_F2_50 ,
 REGofMAX1DataOut_F2_52 , REGofMAX1DataOut_F2_54 , REGofMAX1DataOut_F2_56 , REGofMAX1DataOut_F2_58 , REGofMAX1DataOut_F2_74 , REGofMAX1DataOut_F2_76 ,REGofMAX1DataOut_F2_78  ,
 REGofMAX1DataOut_F2_80, REGofMAX1DataOut_F2_82 , REGofMAX1DataOut_F2_98 , REGofMAX1DataOut_F2_100 , REGofMAX1DataOut_F2_102 , REGofMAX1DataOut_F2_104 , REGofMAX1DataOut_F2_106 ,
 REGofMAX1DataOut_F2_122, REGofMAX1DataOut_F2_124 , REGofMAX1DataOut_F2_126 , REGofMAX1DataOut_F2_128 , REGofMAX1DataOut_F2_130 , bigaddress222, Super_2_3_2_1_ch2 );
SUPERMUXMODULECONV2_new mux3_1_2_1_ch2 ( REGofMAX1DataOut_F2_36, REGofMAX1DataOut_F2_38 , REGofMAX1DataOut_F2_40 , REGofMAX1DataOut_F2_42 , REGofMAX1DataOut_F2_44 , REGofMAX1DataOut_F2_60 ,
 REGofMAX1DataOut_F2_62 , REGofMAX1DataOut_F2_64 , REGofMAX1DataOut_F2_66 , REGofMAX1DataOut_F2_68 , REGofMAX1DataOut_F2_84 , REGofMAX1DataOut_F2_86 ,REGofMAX1DataOut_F2_88  ,
 REGofMAX1DataOut_F2_90, REGofMAX1DataOut_F2_92 , REGofMAX1DataOut_F2_108 , REGofMAX1DataOut_F2_110 , REGofMAX1DataOut_F2_112 , REGofMAX1DataOut_F2_114 , REGofMAX1DataOut_F2_116 ,
 REGofMAX1DataOut_F2_132, REGofMAX1DataOut_F2_134 , REGofMAX1DataOut_F2_136 , REGofMAX1DataOut_F2_138 , REGofMAX1DataOut_F2_140 , bigaddress222, Super_3_1_2_1_ch2 );
SUPERMUXMODULECONV2_new mux3_2_2_1_ch2 ( REGofMAX1DataOut_F2_37, REGofMAX1DataOut_F2_39 , REGofMAX1DataOut_F2_41 , REGofMAX1DataOut_F2_43 , REGofMAX1DataOut_F2_45 , REGofMAX1DataOut_F2_61 ,
 REGofMAX1DataOut_F2_63 , REGofMAX1DataOut_F2_65 , REGofMAX1DataOut_F2_67 , REGofMAX1DataOut_F2_69 , REGofMAX1DataOut_F2_85 , REGofMAX1DataOut_F2_87 , REGofMAX1DataOut_F2_89 ,
 REGofMAX1DataOut_F2_91, REGofMAX1DataOut_F2_93 , REGofMAX1DataOut_F2_109 , REGofMAX1DataOut_F2_111 , REGofMAX1DataOut_F2_113 , REGofMAX1DataOut_F2_115 , REGofMAX1DataOut_F2_117 ,
 REGofMAX1DataOut_F2_133, REGofMAX1DataOut_F2_135 , REGofMAX1DataOut_F2_137 , REGofMAX1DataOut_F2_139 , REGofMAX1DataOut_F2_141 , bigaddress222, Super_3_2_2_1_ch2 );
SUPERMUXMODULECONV2_new mux3_3_2_1_ch2 ( REGofMAX1DataOut_F2_38, REGofMAX1DataOut_F2_40 , REGofMAX1DataOut_F2_42 , REGofMAX1DataOut_F2_44 , REGofMAX1DataOut_F2_46 , REGofMAX1DataOut_F2_62 ,
 REGofMAX1DataOut_F2_64 , REGofMAX1DataOut_F2_66 , REGofMAX1DataOut_F2_68 , REGofMAX1DataOut_F2_70 , REGofMAX1DataOut_F2_86 , REGofMAX1DataOut_F2_88 , REGofMAX1DataOut_F2_90 ,
 REGofMAX1DataOut_F2_92, REGofMAX1DataOut_F2_94 , REGofMAX1DataOut_F2_110 , REGofMAX1DataOut_F2_112 , REGofMAX1DataOut_F2_114 , REGofMAX1DataOut_F2_116 , REGofMAX1DataOut_F2_118 ,
 REGofMAX1DataOut_F2_134,  REGofMAX1DataOut_F2_136, REGofMAX1DataOut_F2_138 , REGofMAX1DataOut_F2_140 , REGofMAX1DataOut_F2_142 , bigaddress222, Super_3_3_2_1_ch2 );


SUPERMUXMODULECONV2_new mux1_1_2_2_ch2 ( REGofMAX1DataOut_F2_13, REGofMAX1DataOut_F2_15 , REGofMAX1DataOut_F2_17 , REGofMAX1DataOut_F2_19 , REGofMAX1DataOut_F2_21 , REGofMAX1DataOut_F2_37 ,
 REGofMAX1DataOut_F2_39 , REGofMAX1DataOut_F2_41 , REGofMAX1DataOut_F2_43 , REGofMAX1DataOut_F2_45 , REGofMAX1DataOut_F2_61 , REGofMAX1DataOut_F2_63 , REGofMAX1DataOut_F2_65 ,
 REGofMAX1DataOut_F2_67, REGofMAX1DataOut_F2_69 , REGofMAX1DataOut_F2_85 , REGofMAX1DataOut_F2_87 , REGofMAX1DataOut_F2_89 , REGofMAX1DataOut_F2_91 , REGofMAX1DataOut_F2_93 ,
 REGofMAX1DataOut_F2_109, REGofMAX1DataOut_F2_111 , REGofMAX1DataOut_F2_113 , REGofMAX1DataOut_F2_115 , REGofMAX1DataOut_F2_117 , bigaddress222, Super_1_1_2_2_ch2 );
SUPERMUXMODULECONV2_new mux1_2_2_2_ch2 ( REGofMAX1DataOut_F2_14, REGofMAX1DataOut_F2_16 , REGofMAX1DataOut_F2_18 , REGofMAX1DataOut_F2_20 , REGofMAX1DataOut_F2_22 , REGofMAX1DataOut_F2_38 ,
 REGofMAX1DataOut_F2_40 , REGofMAX1DataOut_F2_42 , REGofMAX1DataOut_F2_44 , REGofMAX1DataOut_F2_46 , REGofMAX1DataOut_F2_62 , REGofMAX1DataOut_F2_64 , REGofMAX1DataOut_F2_66 ,
REGofMAX1DataOut_F2_68 , REGofMAX1DataOut_F2_70 , REGofMAX1DataOut_F2_86 , REGofMAX1DataOut_F2_88 , REGofMAX1DataOut_F2_90 , REGofMAX1DataOut_F2_92 , REGofMAX1DataOut_F2_94 ,
 REGofMAX1DataOut_F2_110 , REGofMAX1DataOut_F2_112 , REGofMAX1DataOut_F2_114 , REGofMAX1DataOut_F2_116 , REGofMAX1DataOut_F2_118 , bigaddress222, Super_1_2_2_2_ch2 );
SUPERMUXMODULECONV2_new mux1_3_2_2_ch2 ( REGofMAX1DataOut_F2_15, REGofMAX1DataOut_F2_17 , REGofMAX1DataOut_F2_19 , REGofMAX1DataOut_F2_21 , REGofMAX1DataOut_F2_23 , REGofMAX1DataOut_F2_39 ,
 REGofMAX1DataOut_F2_41 , REGofMAX1DataOut_F2_43 , REGofMAX1DataOut_F2_45 , REGofMAX1DataOut_F2_47 , REGofMAX1DataOut_F2_63 , REGofMAX1DataOut_F2_65 , REGofMAX1DataOut_F2_67 ,
 REGofMAX1DataOut_F2_69, REGofMAX1DataOut_F2_71 , REGofMAX1DataOut_F2_87 , REGofMAX1DataOut_F2_89 , REGofMAX1DataOut_F2_91 , REGofMAX1DataOut_F2_93 , REGofMAX1DataOut_F2_95 ,
 REGofMAX1DataOut_F2_111, REGofMAX1DataOut_F2_113 , REGofMAX1DataOut_F2_115 , REGofMAX1DataOut_F2_117 , REGofMAX1DataOut_F2_119 , bigaddress222, Super_1_3_2_2_ch2 );
SUPERMUXMODULECONV2_new mux2_1_2_2_ch2 ( REGofMAX1DataOut_F2_25, REGofMAX1DataOut_F2_27 , REGofMAX1DataOut_F2_29 , REGofMAX1DataOut_F2_31 , REGofMAX1DataOut_F2_33 , REGofMAX1DataOut_F2_49 ,
 REGofMAX1DataOut_F2_51 , REGofMAX1DataOut_F2_53 , REGofMAX1DataOut_F2_55 , REGofMAX1DataOut_F2_57 , REGofMAX1DataOut_F2_73 , REGofMAX1DataOut_F2_75 , REGofMAX1DataOut_F2_77 ,
 REGofMAX1DataOut_F2_79, REGofMAX1DataOut_F2_81 , REGofMAX1DataOut_F2_97 , REGofMAX1DataOut_F2_99 , REGofMAX1DataOut_F2_101 , REGofMAX1DataOut_F2_103 , REGofMAX1DataOut_F2_105 ,
 REGofMAX1DataOut_F2_121, REGofMAX1DataOut_F2_123 , REGofMAX1DataOut_F2_125 , REGofMAX1DataOut_F2_127 , REGofMAX1DataOut_F2_129 , bigaddress222, Super_2_1_2_2_ch2 );
SUPERMUXMODULECONV2_new mux2_2_2_2_ch2 ( REGofMAX1DataOut_F2_26, REGofMAX1DataOut_F2_28 , REGofMAX1DataOut_F2_30 , REGofMAX1DataOut_F2_32 , REGofMAX1DataOut_F2_34 , REGofMAX1DataOut_F2_50 ,
 REGofMAX1DataOut_F2_52 , REGofMAX1DataOut_F2_54 , REGofMAX1DataOut_F2_56 , REGofMAX1DataOut_F2_58 , REGofMAX1DataOut_F2_74 , REGofMAX1DataOut_F2_76 , REGofMAX1DataOut_F2_78 ,
 REGofMAX1DataOut_F2_80, REGofMAX1DataOut_F2_82 , REGofMAX1DataOut_F2_98 , REGofMAX1DataOut_F2_100 , REGofMAX1DataOut_F2_102 , REGofMAX1DataOut_F2_104 , REGofMAX1DataOut_F2_106 ,
 REGofMAX1DataOut_F2_122, REGofMAX1DataOut_F2_124 , REGofMAX1DataOut_F2_126 , REGofMAX1DataOut_F2_128 , REGofMAX1DataOut_F2_130 , bigaddress222, Super_2_2_2_2_ch2 );
SUPERMUXMODULECONV2_new mux2_3_2_2_ch2 ( REGofMAX1DataOut_F2_27, REGofMAX1DataOut_F2_29 , REGofMAX1DataOut_F2_31 , REGofMAX1DataOut_F2_33 , REGofMAX1DataOut_F2_35 , REGofMAX1DataOut_F2_51 ,
 REGofMAX1DataOut_F2_53 , REGofMAX1DataOut_F2_55 , REGofMAX1DataOut_F2_57 , REGofMAX1DataOut_F2_59 , REGofMAX1DataOut_F2_75 , REGofMAX1DataOut_F2_77 , REGofMAX1DataOut_F2_79 ,
 REGofMAX1DataOut_F2_81, REGofMAX1DataOut_F2_83 , REGofMAX1DataOut_F2_99 , REGofMAX1DataOut_F2_101 , REGofMAX1DataOut_F2_103 , REGofMAX1DataOut_F2_105 , REGofMAX1DataOut_F2_107 ,
 REGofMAX1DataOut_F2_123, REGofMAX1DataOut_F2_125 , REGofMAX1DataOut_F2_127 , REGofMAX1DataOut_F2_129 , REGofMAX1DataOut_F2_131 , bigaddress222, Super_2_3_2_2_ch2 );
SUPERMUXMODULECONV2_new mux3_1_2_2_ch2 ( REGofMAX1DataOut_F2_37, REGofMAX1DataOut_F2_39 , REGofMAX1DataOut_F2_41 , REGofMAX1DataOut_F2_43 , REGofMAX1DataOut_F2_45 , REGofMAX1DataOut_F2_61 ,
 REGofMAX1DataOut_F2_63 , REGofMAX1DataOut_F2_65 , REGofMAX1DataOut_F2_67 , REGofMAX1DataOut_F2_69 , REGofMAX1DataOut_F2_85 , REGofMAX1DataOut_F2_87 , REGofMAX1DataOut_F2_89 ,
 REGofMAX1DataOut_F2_91, REGofMAX1DataOut_F2_93 , REGofMAX1DataOut_F2_109 , REGofMAX1DataOut_F2_111 , REGofMAX1DataOut_F2_113 , REGofMAX1DataOut_F2_115 , REGofMAX1DataOut_F2_117 ,
 REGofMAX1DataOut_F2_133, REGofMAX1DataOut_F2_135 ,REGofMAX1DataOut_F2_137  , REGofMAX1DataOut_F2_139 , REGofMAX1DataOut_F2_141 , bigaddress222, Super_3_1_2_2_ch2 );
SUPERMUXMODULECONV2_new mux3_2_2_2_ch2 ( REGofMAX1DataOut_F2_38, REGofMAX1DataOut_F2_40 , REGofMAX1DataOut_F2_42 , REGofMAX1DataOut_F2_44 , REGofMAX1DataOut_F2_46 , REGofMAX1DataOut_F2_62 ,
 REGofMAX1DataOut_F2_64 , REGofMAX1DataOut_F2_66 , REGofMAX1DataOut_F2_68 , REGofMAX1DataOut_F2_70 , REGofMAX1DataOut_F2_86 , REGofMAX1DataOut_F2_88 , REGofMAX1DataOut_F2_90 ,
 REGofMAX1DataOut_F2_92, REGofMAX1DataOut_F2_94 , REGofMAX1DataOut_F2_110 , REGofMAX1DataOut_F2_112 , REGofMAX1DataOut_F2_114 , REGofMAX1DataOut_F2_116 , REGofMAX1DataOut_F2_118 ,
REGofMAX1DataOut_F2_134 , REGofMAX1DataOut_F2_136 , REGofMAX1DataOut_F2_138 , REGofMAX1DataOut_F2_140 , REGofMAX1DataOut_F2_142 , bigaddress222, Super_3_2_2_2_ch2 );
SUPERMUXMODULECONV2_new mux3_3_2_2_ch2 ( REGofMAX1DataOut_F2_39, REGofMAX1DataOut_F2_41 , REGofMAX1DataOut_F2_43 , REGofMAX1DataOut_F2_45 , REGofMAX1DataOut_F2_47 , REGofMAX1DataOut_F2_63 ,
 REGofMAX1DataOut_F2_65 , REGofMAX1DataOut_F2_67 , REGofMAX1DataOut_F2_69 , REGofMAX1DataOut_F2_71 , REGofMAX1DataOut_F2_87 , REGofMAX1DataOut_F2_89 , REGofMAX1DataOut_F2_91 ,
 REGofMAX1DataOut_F2_93, REGofMAX1DataOut_F2_95 , REGofMAX1DataOut_F2_111 , REGofMAX1DataOut_F2_113 , REGofMAX1DataOut_F2_115 , REGofMAX1DataOut_F2_117 , REGofMAX1DataOut_F2_119 ,
 REGofMAX1DataOut_F2_135, REGofMAX1DataOut_F2_137 , REGofMAX1DataOut_F2_139 , REGofMAX1DataOut_F2_141 ,  REGofMAX1DataOut_F2_143, bigaddress222, Super_3_3_2_2_ch2 );

MUX9X1_conv2 In2_CONV2_MUX0 ( Super_1_1_1_1_ch2 , Super_1_2_1_1_ch2 , Super_1_3_1_1_ch2 , Super_2_1_1_1_ch2 , Super_2_2_1_1_ch2 , Super_2_3_1_1_ch2 , Super_3_1_1_1_ch2 , Super_3_2_1_1_ch2 , Super_3_3_1_1_ch2  ,  CONV2_address , In2_CONV2_MUXout0 );
MUX9X1_conv2 In2_CONV2_MUX1 ( Super_1_1_1_2_ch2 , Super_1_2_1_2_ch2 , Super_1_3_1_2_ch2 , Super_2_1_1_2_ch2 , Super_2_2_1_2_ch2 , Super_2_3_1_2_ch2 , Super_3_1_1_2_ch2 ,   Super_3_2_1_2_ch2 , Super_3_3_1_2_ch2 ,  CONV2_address , In2_CONV2_MUXout1 );
MUX9X1_conv2 In2_CONV2_MUX10 ( Super_1_1_2_1_ch2 , Super_1_2_2_1_ch2 , Super_1_3_2_1_ch2 , Super_2_1_2_1_ch2 , Super_2_2_2_1_ch2 , Super_2_3_2_1_ch2 , Super_3_1_2_1_ch2 , Super_3_2_2_1_ch2 , Super_3_3_2_1_ch2   ,  CONV2_address , In2_CONV2_MUXout10 );
MUX9X1_conv2 In2_CONV2_MUX11 (  Super_1_1_2_2_ch2 , Super_1_2_2_2_ch2 , Super_1_3_2_2_ch2 , Super_2_1_2_2_ch2 , Super_2_2_2_2_ch2 , Super_2_3_2_2_ch2 , Super_3_1_2_2_ch2 ,  Super_3_2_2_2_ch2 , Super_3_3_2_2_ch2  ,  CONV2_address , In2_CONV2_MUXout11 );





MAC_9 In2_CONV2_MAC0_F1 (In2_CONV2_ROMout, In2_CONV2_MUXout0 , clk, In2_CONV2_MACoutF1_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC1_F1  (In2_CONV2_ROMout, In2_CONV2_MUXout1 , clk, In2_CONV2_MACoutF1_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC10_F1  (In2_CONV2_ROMout, In2_CONV2_MUXout10 , clk, In2_CONV2_MACoutF1_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC11_F1  (In2_CONV2_ROMout, In2_CONV2_MUXout11 , clk, In2_CONV2_MACoutF1_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In2_CONV2_MAC0_F2 (In2_CONV2_ROMout1, In2_CONV2_MUXout0 , clk, In2_CONV2_MACoutF2_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC1_F2  (In2_CONV2_ROMout1, In2_CONV2_MUXout1 , clk, In2_CONV2_MACoutF2_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC10_F2  (In2_CONV2_ROMout1, In2_CONV2_MUXout10 , clk, In2_CONV2_MACoutF2_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC11_F2  (In2_CONV2_ROMout1, In2_CONV2_MUXout11 , clk, In2_CONV2_MACoutF2_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In2_CONV2_MAC0_F3 (In2_CONV2_ROMout2, In2_CONV2_MUXout0 , clk, In2_CONV2_MACoutF3_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC1_F3 (In2_CONV2_ROMout2, In2_CONV2_MUXout1 , clk, In2_CONV2_MACoutF3_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC10_F3 (In2_CONV2_ROMout2, In2_CONV2_MUXout10 , clk, In2_CONV2_MACoutF3_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC11_F3 (In2_CONV2_ROMout2, In2_CONV2_MUXout11 , clk, In2_CONV2_MACoutF3_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In2_CONV2_MAC0_F4 (In2_CONV2_ROMout3, In2_CONV2_MUXout0 , clk, In2_CONV2_MACoutF4_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC1_F4  (In2_CONV2_ROMout3, In2_CONV2_MUXout1 , clk, In2_CONV2_MACoutF4_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC10_F4  (In2_CONV2_ROMout3, In2_CONV2_MUXout10 , clk, In2_CONV2_MACoutF4_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In2_CONV2_MAC11_F4  (In2_CONV2_ROMout3, In2_CONV2_MUXout11 , clk, In2_CONV2_MACoutF4_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

//3rd input

SUPERMUXMODULECONV2_new mux1_1_1_1_ch3 ( REGofMAX1DataOut_F3_0, REGofMAX1DataOut_F3_2 , REGofMAX1DataOut_F3_4 , REGofMAX1DataOut_F3_6 , REGofMAX1DataOut_F3_8 , REGofMAX1DataOut_F3_24 ,
 REGofMAX1DataOut_F3_26 , REGofMAX1DataOut_F3_28 , REGofMAX1DataOut_F3_30 , REGofMAX1DataOut_F3_32 , REGofMAX1DataOut_F3_48 , REGofMAX1DataOut_F3_50 , REGofMAX1DataOut_F3_52 ,
 REGofMAX1DataOut_F3_54, REGofMAX1DataOut_F3_56 , REGofMAX1DataOut_F3_72 , REGofMAX1DataOut_F3_74 , REGofMAX1DataOut_F3_76 , REGofMAX1DataOut_F3_78 , REGofMAX1DataOut_F3_80 ,
 REGofMAX1DataOut_F3_96, REGofMAX1DataOut_F3_98 ,REGofMAX1DataOut_F3_100  , REGofMAX1DataOut_F3_102 , REGofMAX1DataOut_F3_104 , bigaddress222, Super_1_1_1_1_ch3 );
SUPERMUXMODULECONV2_new mux1_2_1_1_ch3 ( REGofMAX1DataOut_F3_1 , REGofMAX1DataOut_F3_3 , REGofMAX1DataOut_F3_5 , REGofMAX1DataOut_F3_7 , REGofMAX1DataOut_F3_9 , REGofMAX1DataOut_F3_25 ,
 REGofMAX1DataOut_F3_27 , REGofMAX1DataOut_F3_29 , REGofMAX1DataOut_F3_31 , REGofMAX1DataOut_F3_33 , REGofMAX1DataOut_F3_49 , REGofMAX1DataOut_F3_51 , REGofMAX1DataOut_F3_53 ,
 REGofMAX1DataOut_F3_55, REGofMAX1DataOut_F3_57 , REGofMAX1DataOut_F3_73 , REGofMAX1DataOut_F3_75 , REGofMAX1DataOut_F3_77 , REGofMAX1DataOut_F3_79 , REGofMAX1DataOut_F3_81 ,
 REGofMAX1DataOut_F3_97, REGofMAX1DataOut_F3_99 , REGofMAX1DataOut_F3_101 , REGofMAX1DataOut_F3_103 ,  REGofMAX1DataOut_F3_105, bigaddress222, Super_1_2_1_1_ch3 );
SUPERMUXMODULECONV2_new mux1_3_1_1_ch3 ( REGofMAX1DataOut_F3_2,  REGofMAX1DataOut_F3_4, REGofMAX1DataOut_F3_6 , REGofMAX1DataOut_F3_8 , REGofMAX1DataOut_F3_10 , REGofMAX1DataOut_F3_26 ,
 REGofMAX1DataOut_F3_28 , REGofMAX1DataOut_F3_30 , REGofMAX1DataOut_F3_32 , REGofMAX1DataOut_F3_34 , REGofMAX1DataOut_F3_50 , REGofMAX1DataOut_F3_52 , REGofMAX1DataOut_F3_54 ,
 REGofMAX1DataOut_F3_56, REGofMAX1DataOut_F3_58 , REGofMAX1DataOut_F3_74 , REGofMAX1DataOut_F3_76 , REGofMAX1DataOut_F3_78 , REGofMAX1DataOut_F3_80 , REGofMAX1DataOut_F3_82 ,
 REGofMAX1DataOut_F3_98, REGofMAX1DataOut_F3_100 , REGofMAX1DataOut_F3_102 , REGofMAX1DataOut_F3_104 , REGofMAX1DataOut_F3_106 , bigaddress222, Super_1_3_1_1_ch3 );
SUPERMUXMODULECONV2_new mux2_1_1_1_ch3 ( REGofMAX1DataOut_F3_12 ,REGofMAX1DataOut_F3_14  , REGofMAX1DataOut_F3_16 , REGofMAX1DataOut_F3_18 , REGofMAX1DataOut_F3_20 , REGofMAX1DataOut_F3_36 ,
 REGofMAX1DataOut_F3_38 , REGofMAX1DataOut_F3_40 , REGofMAX1DataOut_F3_42 , REGofMAX1DataOut_F3_44 , REGofMAX1DataOut_F3_60 , REGofMAX1DataOut_F3_62 , REGofMAX1DataOut_F3_64 ,
 REGofMAX1DataOut_F3_66, REGofMAX1DataOut_F3_68 , REGofMAX1DataOut_F3_84 , REGofMAX1DataOut_F3_86 , REGofMAX1DataOut_F3_88 , REGofMAX1DataOut_F3_90 , REGofMAX1DataOut_F3_92  ,
 REGofMAX1DataOut_F3_108, REGofMAX1DataOut_F3_110 , REGofMAX1DataOut_F3_112 , REGofMAX1DataOut_F3_114 , REGofMAX1DataOut_F3_116 , bigaddress222, Super_2_1_1_1_ch3 );
SUPERMUXMODULECONV2_new mux2_2_1_1_ch3 ( REGofMAX1DataOut_F3_13, REGofMAX1DataOut_F3_15 , REGofMAX1DataOut_F3_17 , REGofMAX1DataOut_F3_19 , REGofMAX1DataOut_F3_21 , REGofMAX1DataOut_F3_37 ,
 REGofMAX1DataOut_F3_39 , REGofMAX1DataOut_F3_41 , REGofMAX1DataOut_F3_43 , REGofMAX1DataOut_F3_45 , REGofMAX1DataOut_F3_61 , REGofMAX1DataOut_F3_63 , REGofMAX1DataOut_F3_65 ,
 REGofMAX1DataOut_F3_67, REGofMAX1DataOut_F3_69 , REGofMAX1DataOut_F3_85 , REGofMAX1DataOut_F3_87 , REGofMAX1DataOut_F3_89 , REGofMAX1DataOut_F3_91 ,REGofMAX1DataOut_F3_93  ,
 REGofMAX1DataOut_F3_109, REGofMAX1DataOut_F3_111 , REGofMAX1DataOut_F3_113 , REGofMAX1DataOut_F3_115 ,REGofMAX1DataOut_F3_117  , bigaddress222, Super_2_2_1_1_ch3 );
SUPERMUXMODULECONV2_new mux2_3_1_1_ch3 ( REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_16  , REGofMAX1DataOut_F3_18 , REGofMAX1DataOut_F3_20 , REGofMAX1DataOut_F3_22 , REGofMAX1DataOut_F3_38 ,
 REGofMAX1DataOut_F3_40 , REGofMAX1DataOut_F3_42 , REGofMAX1DataOut_F3_44 , REGofMAX1DataOut_F3_46 , REGofMAX1DataOut_F3_62 , REGofMAX1DataOut_F3_64 , REGofMAX1DataOut_F3_66 ,
 REGofMAX1DataOut_F3_68, REGofMAX1DataOut_F3_70 , REGofMAX1DataOut_F3_86 , REGofMAX1DataOut_F3_88 , REGofMAX1DataOut_F3_90 , REGofMAX1DataOut_F3_92 , REGofMAX1DataOut_F3_94 ,
 REGofMAX1DataOut_F3_110, REGofMAX1DataOut_F3_112 , REGofMAX1DataOut_F3_114 , REGofMAX1DataOut_F3_116 , REGofMAX1DataOut_F3_118 , bigaddress222, Super_2_3_1_1_ch3 );
SUPERMUXMODULECONV2_new mux3_1_1_1_ch3 ( REGofMAX1DataOut_F3_24, REGofMAX1DataOut_F3_26 , REGofMAX1DataOut_F3_28 , REGofMAX1DataOut_F3_30 , REGofMAX1DataOut_F3_32 , REGofMAX1DataOut_F3_48 ,
 REGofMAX1DataOut_F3_50 , REGofMAX1DataOut_F3_52 , REGofMAX1DataOut_F3_54 , REGofMAX1DataOut_F3_56 , REGofMAX1DataOut_F3_72 , REGofMAX1DataOut_F3_74 , REGofMAX1DataOut_F3_76 ,
 REGofMAX1DataOut_F3_78, REGofMAX1DataOut_F3_80 , REGofMAX1DataOut_F3_96 , REGofMAX1DataOut_F3_98 , REGofMAX1DataOut_F3_100 , REGofMAX1DataOut_F3_102 , REGofMAX1DataOut_F3_104 ,
 REGofMAX1DataOut_F3_120, REGofMAX1DataOut_F3_122 , REGofMAX1DataOut_F3_124 , REGofMAX1DataOut_F3_126 , REGofMAX1DataOut_F3_128 , bigaddress222, Super_3_1_1_1_ch3 );
SUPERMUXMODULECONV2_new mux3_2_1_1_ch3 ( REGofMAX1DataOut_F3_25, REGofMAX1DataOut_F3_27 , REGofMAX1DataOut_F3_29 , REGofMAX1DataOut_F3_31 , REGofMAX1DataOut_F3_33 , REGofMAX1DataOut_F3_49 ,
 REGofMAX1DataOut_F3_51 ,REGofMAX1DataOut_F3_53  , REGofMAX1DataOut_F3_55 , REGofMAX1DataOut_F3_57 , REGofMAX1DataOut_F3_73 , REGofMAX1DataOut_F3_75 , REGofMAX1DataOut_F3_77 ,
REGofMAX1DataOut_F3_79 , REGofMAX1DataOut_F3_81 , REGofMAX1DataOut_F3_97 , REGofMAX1DataOut_F3_99 , REGofMAX1DataOut_F3_101 , REGofMAX1DataOut_F3_103 , REGofMAX1DataOut_F3_105 ,
 REGofMAX1DataOut_F3_121 , REGofMAX1DataOut_F3_123 , REGofMAX1DataOut_F3_125 , REGofMAX1DataOut_F3_127 , REGofMAX1DataOut_F3_129 , bigaddress222, Super_3_2_1_1_ch3 );
SUPERMUXMODULECONV2_new mux3_3_1_1_ch3 ( REGofMAX1DataOut_F3_26, REGofMAX1DataOut_F3_28 , REGofMAX1DataOut_F3_30 , REGofMAX1DataOut_F3_32 , REGofMAX1DataOut_F3_34 , REGofMAX1DataOut_F3_50 ,
REGofMAX1DataOut_F3_52  , REGofMAX1DataOut_F3_54 , REGofMAX1DataOut_F3_56 , REGofMAX1DataOut_F3_58 , REGofMAX1DataOut_F3_74 , REGofMAX1DataOut_F3_76 , REGofMAX1DataOut_F3_78 ,
REGofMAX1DataOut_F3_80 , REGofMAX1DataOut_F3_82 , REGofMAX1DataOut_F3_98 , REGofMAX1DataOut_F3_100 , REGofMAX1DataOut_F3_102 , REGofMAX1DataOut_F3_104 , REGofMAX1DataOut_F3_106 ,
 REGofMAX1DataOut_F3_122 , REGofMAX1DataOut_F3_124 , REGofMAX1DataOut_F3_126 , REGofMAX1DataOut_F3_128 , REGofMAX1DataOut_F3_130 , bigaddress222, Super_3_3_1_1_ch3 );



SUPERMUXMODULECONV2_new mux1_1_1_2_ch3 ( REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_3  , REGofMAX1DataOut_F3_5 , REGofMAX1DataOut_F3_7 , REGofMAX1DataOut_F3_9 , REGofMAX1DataOut_F3_25 ,
REGofMAX1DataOut_F3_27 , REGofMAX1DataOut_F3_29 , REGofMAX1DataOut_F3_31 , REGofMAX1DataOut_F3_33 , REGofMAX1DataOut_F3_49 , REGofMAX1DataOut_F3_51 ,REGofMAX1DataOut_F3_53  ,
 REGofMAX1DataOut_F3_55 ,REGofMAX1DataOut_F3_57  , REGofMAX1DataOut_F3_73 , REGofMAX1DataOut_F3_75 , REGofMAX1DataOut_F3_77 , REGofMAX1DataOut_F3_79 , REGofMAX1DataOut_F3_81 ,
 REGofMAX1DataOut_F3_97, REGofMAX1DataOut_F3_99 , REGofMAX1DataOut_F3_101 , REGofMAX1DataOut_F3_103 , REGofMAX1DataOut_F3_105 , bigaddress222, Super_1_1_1_2_ch3 );
SUPERMUXMODULECONV2_new mux1_2_1_2_ch3 ( REGofMAX1DataOut_F3_2, REGofMAX1DataOut_F3_4 , REGofMAX1DataOut_F3_6 , REGofMAX1DataOut_F3_8 , REGofMAX1DataOut_F3_10 , REGofMAX1DataOut_F3_26 ,
REGofMAX1DataOut_F3_28 , REGofMAX1DataOut_F3_30 , REGofMAX1DataOut_F3_32 , REGofMAX1DataOut_F3_34 , REGofMAX1DataOut_F3_50 , REGofMAX1DataOut_F3_52 ,REGofMAX1DataOut_F3_54  ,
 REGofMAX1DataOut_F3_56 , REGofMAX1DataOut_F3_58 , REGofMAX1DataOut_F3_74 , REGofMAX1DataOut_F3_76 , REGofMAX1DataOut_F3_78 , REGofMAX1DataOut_F3_80 , REGofMAX1DataOut_F3_82 ,
 REGofMAX1DataOut_F3_98, REGofMAX1DataOut_F3_100 , REGofMAX1DataOut_F3_102 , REGofMAX1DataOut_F3_104 , REGofMAX1DataOut_F3_106 , bigaddress222, Super_1_2_1_2_ch3 );
SUPERMUXMODULECONV2_new mux1_3_1_2_ch3 ( REGofMAX1DataOut_F3_3, REGofMAX1DataOut_F3_5 , REGofMAX1DataOut_F3_7 , REGofMAX1DataOut_F3_9 , REGofMAX1DataOut_F3_11 , REGofMAX1DataOut_F3_27 ,
REGofMAX1DataOut_F3_29 , REGofMAX1DataOut_F3_31 , REGofMAX1DataOut_F3_33 , REGofMAX1DataOut_F3_35 , REGofMAX1DataOut_F3_51 , REGofMAX1DataOut_F3_53 , REGofMAX1DataOut_F3_55 ,
 REGofMAX1DataOut_F3_57 , REGofMAX1DataOut_F3_59 , REGofMAX1DataOut_F3_75 , REGofMAX1DataOut_F3_77 , REGofMAX1DataOut_F3_79 , REGofMAX1DataOut_F3_81 , REGofMAX1DataOut_F3_83 ,
 REGofMAX1DataOut_F3_99, REGofMAX1DataOut_F3_101 , REGofMAX1DataOut_F3_103 , REGofMAX1DataOut_F3_105 , REGofMAX1DataOut_F3_107 , bigaddress222, Super_1_3_1_2_ch3 );
SUPERMUXMODULECONV2_new mux2_1_1_2_ch3 ( REGofMAX1DataOut_F3_13, REGofMAX1DataOut_F3_15 , REGofMAX1DataOut_F3_17 , REGofMAX1DataOut_F3_19 , REGofMAX1DataOut_F3_21 , REGofMAX1DataOut_F3_37 ,
REGofMAX1DataOut_F3_39 , REGofMAX1DataOut_F3_41 , REGofMAX1DataOut_F3_43 , REGofMAX1DataOut_F3_45 , REGofMAX1DataOut_F3_61 , REGofMAX1DataOut_F3_63  ,REGofMAX1DataOut_F3_65  ,
 REGofMAX1DataOut_F3_67 , REGofMAX1DataOut_F3_69 , REGofMAX1DataOut_F3_85 , REGofMAX1DataOut_F3_87 , REGofMAX1DataOut_F3_89 , REGofMAX1DataOut_F3_91 , REGofMAX1DataOut_F3_93 ,
 REGofMAX1DataOut_F3_109, REGofMAX1DataOut_F3_111 , REGofMAX1DataOut_F3_113 , REGofMAX1DataOut_F3_115 , REGofMAX1DataOut_F3_117 , bigaddress222, Super_2_1_1_2_ch3 );
SUPERMUXMODULECONV2_new mux2_2_1_2_ch3 ( REGofMAX1DataOut_F3_14, REGofMAX1DataOut_F3_16 , REGofMAX1DataOut_F3_18 , REGofMAX1DataOut_F3_20 , REGofMAX1DataOut_F3_22 , REGofMAX1DataOut_F3_38 ,
REGofMAX1DataOut_F3_40  , REGofMAX1DataOut_F3_42 , REGofMAX1DataOut_F3_44 , REGofMAX1DataOut_F3_46 , REGofMAX1DataOut_F3_62 , REGofMAX1DataOut_F3_64 ,REGofMAX1DataOut_F3_66  ,
 REGofMAX1DataOut_F3_68 , REGofMAX1DataOut_F3_70 , REGofMAX1DataOut_F3_86 , REGofMAX1DataOut_F3_88 , REGofMAX1DataOut_F3_90 , REGofMAX1DataOut_F3_92 , REGofMAX1DataOut_F3_94 ,
 REGofMAX1DataOut_F3_110, REGofMAX1DataOut_F3_112 , REGofMAX1DataOut_F3_114 , REGofMAX1DataOut_F3_116 , REGofMAX1DataOut_F3_118 , bigaddress222, Super_2_2_1_2_ch3 );
SUPERMUXMODULECONV2_new mux2_3_1_2_ch3 ( REGofMAX1DataOut_F3_15, REGofMAX1DataOut_F3_17 , REGofMAX1DataOut_F3_19 , REGofMAX1DataOut_F3_21 , REGofMAX1DataOut_F3_23 , REGofMAX1DataOut_F3_39 ,
REGofMAX1DataOut_F3_41  , REGofMAX1DataOut_F3_43 , REGofMAX1DataOut_F3_45 , REGofMAX1DataOut_F3_47 , REGofMAX1DataOut_F3_63 , REGofMAX1DataOut_F3_65 ,REGofMAX1DataOut_F3_67  ,
 REGofMAX1DataOut_F3_69 , REGofMAX1DataOut_F3_71 , REGofMAX1DataOut_F3_87 , REGofMAX1DataOut_F3_89 , REGofMAX1DataOut_F3_91 , REGofMAX1DataOut_F3_93 , REGofMAX1DataOut_F3_95 ,
 REGofMAX1DataOut_F3_111, REGofMAX1DataOut_F3_113 , REGofMAX1DataOut_F3_115 , REGofMAX1DataOut_F3_117 , REGofMAX1DataOut_F3_119 , bigaddress222, Super_2_3_1_2_ch3 );
SUPERMUXMODULECONV2_new mux3_1_1_2_ch3 ( REGofMAX1DataOut_F3_25, REGofMAX1DataOut_F3_27 , REGofMAX1DataOut_F3_29 , REGofMAX1DataOut_F3_31 , REGofMAX1DataOut_F3_33 , REGofMAX1DataOut_F3_49 ,
REGofMAX1DataOut_F3_51 , REGofMAX1DataOut_F3_53 , REGofMAX1DataOut_F3_55 , REGofMAX1DataOut_F3_57 , REGofMAX1DataOut_F3_73 , REGofMAX1DataOut_F3_75 ,REGofMAX1DataOut_F3_77  ,
 REGofMAX1DataOut_F3_79 , REGofMAX1DataOut_F3_81 , REGofMAX1DataOut_F3_97 , REGofMAX1DataOut_F3_99 , REGofMAX1DataOut_F3_101 , REGofMAX1DataOut_F3_103 , REGofMAX1DataOut_F3_105 ,
REGofMAX1DataOut_F3_121 , REGofMAX1DataOut_F3_123 , REGofMAX1DataOut_F3_125 , REGofMAX1DataOut_F3_127 , REGofMAX1DataOut_F3_129 , bigaddress222, Super_3_1_1_2_ch3 );
SUPERMUXMODULECONV2_new mux3_2_1_2_ch3 ( REGofMAX1DataOut_F3_26, REGofMAX1DataOut_F3_28 , REGofMAX1DataOut_F3_30 , REGofMAX1DataOut_F3_32 , REGofMAX1DataOut_F3_34 , REGofMAX1DataOut_F3_50 ,
REGofMAX1DataOut_F3_52  , REGofMAX1DataOut_F3_54 , REGofMAX1DataOut_F3_56 , REGofMAX1DataOut_F3_58 , REGofMAX1DataOut_F3_74 , REGofMAX1DataOut_F3_76 ,REGofMAX1DataOut_F3_78  ,
 REGofMAX1DataOut_F3_80 , REGofMAX1DataOut_F3_82 , REGofMAX1DataOut_F3_98 , REGofMAX1DataOut_F3_100 , REGofMAX1DataOut_F3_102 , REGofMAX1DataOut_F3_104 ,REGofMAX1DataOut_F3_106  ,
 REGofMAX1DataOut_F3_122, REGofMAX1DataOut_F3_124 , REGofMAX1DataOut_F3_126 , REGofMAX1DataOut_F3_128 , REGofMAX1DataOut_F3_130 , bigaddress222, Super_3_2_1_2_ch3 );
SUPERMUXMODULECONV2_new mux3_3_1_2_ch3 ( REGofMAX1DataOut_F3_27, REGofMAX1DataOut_F3_29 , REGofMAX1DataOut_F3_31 , REGofMAX1DataOut_F3_33 , REGofMAX1DataOut_F3_35 , REGofMAX1DataOut_F3_51 ,
REGofMAX1DataOut_F3_53 , REGofMAX1DataOut_F3_55 , REGofMAX1DataOut_F3_57 , REGofMAX1DataOut_F3_59 , REGofMAX1DataOut_F3_75 , REGofMAX1DataOut_F3_77 , REGofMAX1DataOut_F3_79 ,
 REGofMAX1DataOut_F3_81 , REGofMAX1DataOut_F3_83 ,REGofMAX1DataOut_F3_99  , REGofMAX1DataOut_F3_101 , REGofMAX1DataOut_F3_103 , REGofMAX1DataOut_F3_105 , REGofMAX1DataOut_F3_107 ,
 REGofMAX1DataOut_F3_123, REGofMAX1DataOut_F3_125 , REGofMAX1DataOut_F3_127 , REGofMAX1DataOut_F3_129 , REGofMAX1DataOut_F3_131 , bigaddress222, Super_3_3_1_2_ch3 );


SUPERMUXMODULECONV2_new mux1_1_2_1_ch3 ( REGofMAX1DataOut_F3_12, REGofMAX1DataOut_F3_14 , REGofMAX1DataOut_F3_16 , REGofMAX1DataOut_F3_18 , REGofMAX1DataOut_F3_20 , REGofMAX1DataOut_F3_36 ,
 REGofMAX1DataOut_F3_38 , REGofMAX1DataOut_F3_40 , REGofMAX1DataOut_F3_42 , REGofMAX1DataOut_F3_44 , REGofMAX1DataOut_F3_60 , REGofMAX1DataOut_F3_62 , REGofMAX1DataOut_F3_64 ,
 REGofMAX1DataOut_F3_66, REGofMAX1DataOut_F3_68 , REGofMAX1DataOut_F3_84 , REGofMAX1DataOut_F3_86 , REGofMAX1DataOut_F3_88 , REGofMAX1DataOut_F3_90 , REGofMAX1DataOut_F3_92 ,
 REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_110  , REGofMAX1DataOut_F3_112 , REGofMAX1DataOut_F3_114 , REGofMAX1DataOut_F3_116 , bigaddress222, Super_1_1_2_1_ch3 );
SUPERMUXMODULECONV2_new mux1_2_2_1_ch3 ( REGofMAX1DataOut_F3_13, REGofMAX1DataOut_F3_15 , REGofMAX1DataOut_F3_17 , REGofMAX1DataOut_F3_19 , REGofMAX1DataOut_F3_21 , REGofMAX1DataOut_F3_37 ,
 REGofMAX1DataOut_F3_39 , REGofMAX1DataOut_F3_41 , REGofMAX1DataOut_F3_43 , REGofMAX1DataOut_F3_45 , REGofMAX1DataOut_F3_61 , REGofMAX1DataOut_F3_63 , REGofMAX1DataOut_F3_65 ,
 REGofMAX1DataOut_F3_67, REGofMAX1DataOut_F3_69 , REGofMAX1DataOut_F3_85 , REGofMAX1DataOut_F3_87 , REGofMAX1DataOut_F3_89 , REGofMAX1DataOut_F3_91 , REGofMAX1DataOut_F3_93 ,
 REGofMAX1DataOut_F3_109, REGofMAX1DataOut_F3_111 , REGofMAX1DataOut_F3_113 , REGofMAX1DataOut_F3_115 , REGofMAX1DataOut_F3_117 , bigaddress222, Super_1_2_2_1_ch3 );
SUPERMUXMODULECONV2_new mux1_3_2_1_ch3 ( REGofMAX1DataOut_F3_14, REGofMAX1DataOut_F3_16 , REGofMAX1DataOut_F3_18 , REGofMAX1DataOut_F3_20 , REGofMAX1DataOut_F3_22 , REGofMAX1DataOut_F3_38 ,
REGofMAX1DataOut_F3_40  , REGofMAX1DataOut_F3_42 , REGofMAX1DataOut_F3_44 , REGofMAX1DataOut_F3_46 , REGofMAX1DataOut_F3_62 , REGofMAX1DataOut_F3_64 ,REGofMAX1DataOut_F3_66 ,
 REGofMAX1DataOut_F3_68 , REGofMAX1DataOut_F3_70 , REGofMAX1DataOut_F3_86 , REGofMAX1DataOut_F3_88 ,REGofMAX1DataOut_F3_90  , REGofMAX1DataOut_F3_92 , REGofMAX1DataOut_F3_94 ,
REGofMAX1DataOut_F3_110 , REGofMAX1DataOut_F3_112 , REGofMAX1DataOut_F3_114 , REGofMAX1DataOut_F3_116 , REGofMAX1DataOut_F3_118 , bigaddress222, Super_1_3_2_1_ch3 );
SUPERMUXMODULECONV2_new mux2_1_2_1_ch3 ( REGofMAX1DataOut_F3_24, REGofMAX1DataOut_F3_26 , REGofMAX1DataOut_F3_28 , REGofMAX1DataOut_F3_30 , REGofMAX1DataOut_F3_32 , REGofMAX1DataOut_F3_48 ,
 REGofMAX1DataOut_F3_50 , REGofMAX1DataOut_F3_52 , REGofMAX1DataOut_F3_54 , REGofMAX1DataOut_F3_56 , REGofMAX1DataOut_F3_72 , REGofMAX1DataOut_F3_74 ,REGofMAX1DataOut_F3_76  ,
 REGofMAX1DataOut_F3_78, REGofMAX1DataOut_F3_80 , REGofMAX1DataOut_F3_96 , REGofMAX1DataOut_F3_98 , REGofMAX1DataOut_F3_100 , REGofMAX1DataOut_F3_102 , REGofMAX1DataOut_F3_104 ,
REGofMAX1DataOut_F3_120 , REGofMAX1DataOut_F3_122 , REGofMAX1DataOut_F3_124 , REGofMAX1DataOut_F3_126 , REGofMAX1DataOut_F3_128 , bigaddress222, Super_2_1_2_1_ch3 );
SUPERMUXMODULECONV2_new mux2_2_2_1_ch3 ( REGofMAX1DataOut_F3_25, REGofMAX1DataOut_F3_27 , REGofMAX1DataOut_F3_29 , REGofMAX1DataOut_F3_31 , REGofMAX1DataOut_F3_33 , REGofMAX1DataOut_F3_49 ,
 REGofMAX1DataOut_F3_51 , REGofMAX1DataOut_F3_53 , REGofMAX1DataOut_F3_55 , REGofMAX1DataOut_F3_57 , REGofMAX1DataOut_F3_73 , REGofMAX1DataOut_F3_75 , REGofMAX1DataOut_F3_77 ,
 REGofMAX1DataOut_F3_79, REGofMAX1DataOut_F3_81 , REGofMAX1DataOut_F3_97 , REGofMAX1DataOut_F3_99 , REGofMAX1DataOut_F3_101 , REGofMAX1DataOut_F3_103 , REGofMAX1DataOut_F3_105 ,
REGofMAX1DataOut_F3_121 , REGofMAX1DataOut_F3_123 , REGofMAX1DataOut_F3_125 , REGofMAX1DataOut_F3_127 , REGofMAX1DataOut_F3_129 , bigaddress222, Super_2_2_2_1_ch3 );
SUPERMUXMODULECONV2_new mux2_3_2_1_ch3 ( REGofMAX1DataOut_F3_26, REGofMAX1DataOut_F3_28 , REGofMAX1DataOut_F3_30 , REGofMAX1DataOut_F3_32 , REGofMAX1DataOut_F3_34 , REGofMAX1DataOut_F3_50 ,
 REGofMAX1DataOut_F3_52 , REGofMAX1DataOut_F3_54 , REGofMAX1DataOut_F3_56 , REGofMAX1DataOut_F3_58 , REGofMAX1DataOut_F3_74 , REGofMAX1DataOut_F3_76 ,REGofMAX1DataOut_F3_78  ,
 REGofMAX1DataOut_F3_80, REGofMAX1DataOut_F3_82 , REGofMAX1DataOut_F3_98 , REGofMAX1DataOut_F3_100 , REGofMAX1DataOut_F3_102 , REGofMAX1DataOut_F3_104 , REGofMAX1DataOut_F3_106 ,
 REGofMAX1DataOut_F3_122, REGofMAX1DataOut_F3_124 , REGofMAX1DataOut_F3_126 , REGofMAX1DataOut_F3_128 , REGofMAX1DataOut_F3_130 , bigaddress222, Super_2_3_2_1_ch3 );
SUPERMUXMODULECONV2_new mux3_1_2_1_ch3 ( REGofMAX1DataOut_F3_36, REGofMAX1DataOut_F3_38 , REGofMAX1DataOut_F3_40 , REGofMAX1DataOut_F3_42 , REGofMAX1DataOut_F3_44 , REGofMAX1DataOut_F3_60 ,
 REGofMAX1DataOut_F3_62 , REGofMAX1DataOut_F3_64 , REGofMAX1DataOut_F3_66 , REGofMAX1DataOut_F3_68 , REGofMAX1DataOut_F3_84 , REGofMAX1DataOut_F3_86 ,REGofMAX1DataOut_F3_88  ,
 REGofMAX1DataOut_F3_90, REGofMAX1DataOut_F3_92 , REGofMAX1DataOut_F3_108 , REGofMAX1DataOut_F3_110 , REGofMAX1DataOut_F3_112 , REGofMAX1DataOut_F3_114 , REGofMAX1DataOut_F3_116 ,
 REGofMAX1DataOut_F3_132, REGofMAX1DataOut_F3_134 , REGofMAX1DataOut_F3_136 , REGofMAX1DataOut_F3_138 , REGofMAX1DataOut_F3_140 , bigaddress222, Super_3_1_2_1_ch3 );
SUPERMUXMODULECONV2_new mux3_2_2_1_ch3 ( REGofMAX1DataOut_F3_37, REGofMAX1DataOut_F3_39 , REGofMAX1DataOut_F3_41 , REGofMAX1DataOut_F3_43 , REGofMAX1DataOut_F3_45 , REGofMAX1DataOut_F3_61 ,
 REGofMAX1DataOut_F3_63 , REGofMAX1DataOut_F3_65 , REGofMAX1DataOut_F3_67 , REGofMAX1DataOut_F3_69 , REGofMAX1DataOut_F3_85 , REGofMAX1DataOut_F3_87 , REGofMAX1DataOut_F3_89 ,
 REGofMAX1DataOut_F3_91, REGofMAX1DataOut_F3_93 , REGofMAX1DataOut_F3_109 , REGofMAX1DataOut_F3_111 , REGofMAX1DataOut_F3_113 , REGofMAX1DataOut_F3_115 , REGofMAX1DataOut_F3_117 ,
 REGofMAX1DataOut_F3_133, REGofMAX1DataOut_F3_135 , REGofMAX1DataOut_F3_137 , REGofMAX1DataOut_F3_139 , REGofMAX1DataOut_F3_141 , bigaddress222, Super_3_2_2_1_ch3 );
SUPERMUXMODULECONV2_new mux3_3_2_1_ch3 ( REGofMAX1DataOut_F3_38, REGofMAX1DataOut_F3_40 , REGofMAX1DataOut_F3_42 , REGofMAX1DataOut_F3_44 , REGofMAX1DataOut_F3_46 , REGofMAX1DataOut_F3_62 ,
 REGofMAX1DataOut_F3_64 , REGofMAX1DataOut_F3_66 , REGofMAX1DataOut_F3_68 , REGofMAX1DataOut_F3_70 , REGofMAX1DataOut_F3_86 , REGofMAX1DataOut_F3_88 , REGofMAX1DataOut_F3_90 ,
 REGofMAX1DataOut_F3_92, REGofMAX1DataOut_F3_94 , REGofMAX1DataOut_F3_110 , REGofMAX1DataOut_F3_112 , REGofMAX1DataOut_F3_114 , REGofMAX1DataOut_F3_116 , REGofMAX1DataOut_F3_118 ,
 REGofMAX1DataOut_F3_134,  REGofMAX1DataOut_F3_136, REGofMAX1DataOut_F3_138 , REGofMAX1DataOut_F3_140 , REGofMAX1DataOut_F3_142 , bigaddress222, Super_3_3_2_1_ch3 );


SUPERMUXMODULECONV2_new mux1_1_2_2_ch3 ( REGofMAX1DataOut_F3_13, REGofMAX1DataOut_F3_15 , REGofMAX1DataOut_F3_17 , REGofMAX1DataOut_F3_19 , REGofMAX1DataOut_F3_21 , REGofMAX1DataOut_F3_37 ,
 REGofMAX1DataOut_F3_39 , REGofMAX1DataOut_F3_41 , REGofMAX1DataOut_F3_43 , REGofMAX1DataOut_F3_45 , REGofMAX1DataOut_F3_61 , REGofMAX1DataOut_F3_63 , REGofMAX1DataOut_F3_65 ,
 REGofMAX1DataOut_F3_67, REGofMAX1DataOut_F3_69 , REGofMAX1DataOut_F3_85 , REGofMAX1DataOut_F3_87 , REGofMAX1DataOut_F3_89 , REGofMAX1DataOut_F3_91 , REGofMAX1DataOut_F3_93 ,
 REGofMAX1DataOut_F3_109, REGofMAX1DataOut_F3_111 , REGofMAX1DataOut_F3_113 , REGofMAX1DataOut_F3_115 , REGofMAX1DataOut_F3_117 , bigaddress222, Super_1_1_2_2_ch3 );
SUPERMUXMODULECONV2_new mux1_2_2_2_ch3 ( REGofMAX1DataOut_F3_14, REGofMAX1DataOut_F3_16 , REGofMAX1DataOut_F3_18 , REGofMAX1DataOut_F3_20 , REGofMAX1DataOut_F3_22 , REGofMAX1DataOut_F3_38 ,
 REGofMAX1DataOut_F3_40 , REGofMAX1DataOut_F3_42 , REGofMAX1DataOut_F3_44 , REGofMAX1DataOut_F3_46 , REGofMAX1DataOut_F3_62 , REGofMAX1DataOut_F3_64 , REGofMAX1DataOut_F3_66 ,
REGofMAX1DataOut_F3_68 , REGofMAX1DataOut_F3_70 , REGofMAX1DataOut_F3_86 , REGofMAX1DataOut_F3_88 , REGofMAX1DataOut_F3_90 , REGofMAX1DataOut_F3_92 , REGofMAX1DataOut_F3_94 ,
 REGofMAX1DataOut_F3_110 , REGofMAX1DataOut_F3_112 , REGofMAX1DataOut_F3_114 , REGofMAX1DataOut_F3_116 , REGofMAX1DataOut_F3_118 , bigaddress222, Super_1_2_2_2_ch3 );
SUPERMUXMODULECONV2_new mux1_3_2_2_ch3 ( REGofMAX1DataOut_F3_15, REGofMAX1DataOut_F3_17 , REGofMAX1DataOut_F3_19 , REGofMAX1DataOut_F3_21 , REGofMAX1DataOut_F3_23 , REGofMAX1DataOut_F3_39 ,
 REGofMAX1DataOut_F3_41 , REGofMAX1DataOut_F3_43 , REGofMAX1DataOut_F3_45 , REGofMAX1DataOut_F3_47 , REGofMAX1DataOut_F3_63 , REGofMAX1DataOut_F3_65 , REGofMAX1DataOut_F3_67 ,
 REGofMAX1DataOut_F3_69, REGofMAX1DataOut_F3_71 , REGofMAX1DataOut_F3_87 , REGofMAX1DataOut_F3_89 , REGofMAX1DataOut_F3_91 , REGofMAX1DataOut_F3_93 , REGofMAX1DataOut_F3_95 ,
 REGofMAX1DataOut_F3_111, REGofMAX1DataOut_F3_113 , REGofMAX1DataOut_F3_115 , REGofMAX1DataOut_F3_117 , REGofMAX1DataOut_F3_119 , bigaddress222, Super_1_3_2_2_ch3 );
SUPERMUXMODULECONV2_new mux2_1_2_2_ch3 ( REGofMAX1DataOut_F3_25, REGofMAX1DataOut_F3_27 , REGofMAX1DataOut_F3_29 , REGofMAX1DataOut_F3_31 , REGofMAX1DataOut_F3_33 , REGofMAX1DataOut_F3_49 ,
 REGofMAX1DataOut_F3_51 , REGofMAX1DataOut_F3_53 , REGofMAX1DataOut_F3_55 , REGofMAX1DataOut_F3_57 , REGofMAX1DataOut_F3_73 , REGofMAX1DataOut_F3_75 , REGofMAX1DataOut_F3_77 ,
 REGofMAX1DataOut_F3_79, REGofMAX1DataOut_F3_81 , REGofMAX1DataOut_F3_97 , REGofMAX1DataOut_F3_99 , REGofMAX1DataOut_F3_101 , REGofMAX1DataOut_F3_103 , REGofMAX1DataOut_F3_105 ,
 REGofMAX1DataOut_F3_121, REGofMAX1DataOut_F3_123 , REGofMAX1DataOut_F3_125 , REGofMAX1DataOut_F3_127 , REGofMAX1DataOut_F3_129 , bigaddress222, Super_2_1_2_2_ch3 );
SUPERMUXMODULECONV2_new mux2_2_2_2_ch3 ( REGofMAX1DataOut_F3_26, REGofMAX1DataOut_F3_28 , REGofMAX1DataOut_F3_30 , REGofMAX1DataOut_F3_32 , REGofMAX1DataOut_F3_34 , REGofMAX1DataOut_F3_50 ,
 REGofMAX1DataOut_F3_52 , REGofMAX1DataOut_F3_54 , REGofMAX1DataOut_F3_56 , REGofMAX1DataOut_F3_58 , REGofMAX1DataOut_F3_74 , REGofMAX1DataOut_F3_76 , REGofMAX1DataOut_F3_78 ,
 REGofMAX1DataOut_F3_80, REGofMAX1DataOut_F3_82 , REGofMAX1DataOut_F3_98 , REGofMAX1DataOut_F3_100 , REGofMAX1DataOut_F3_102 , REGofMAX1DataOut_F3_104 , REGofMAX1DataOut_F3_106 ,
 REGofMAX1DataOut_F3_122, REGofMAX1DataOut_F3_124 , REGofMAX1DataOut_F3_126 , REGofMAX1DataOut_F3_128 , REGofMAX1DataOut_F3_130 , bigaddress222, Super_2_2_2_2_ch3 );
SUPERMUXMODULECONV2_new mux2_3_2_2_ch3 ( REGofMAX1DataOut_F3_27, REGofMAX1DataOut_F3_29 , REGofMAX1DataOut_F3_31 , REGofMAX1DataOut_F3_33 , REGofMAX1DataOut_F3_35 , REGofMAX1DataOut_F3_51 ,
 REGofMAX1DataOut_F3_53 , REGofMAX1DataOut_F3_55 , REGofMAX1DataOut_F3_57 , REGofMAX1DataOut_F3_59 , REGofMAX1DataOut_F3_75 , REGofMAX1DataOut_F3_77 , REGofMAX1DataOut_F3_79 ,
 REGofMAX1DataOut_F3_81, REGofMAX1DataOut_F3_83 , REGofMAX1DataOut_F3_99 , REGofMAX1DataOut_F3_101 , REGofMAX1DataOut_F3_103 , REGofMAX1DataOut_F3_105 , REGofMAX1DataOut_F3_107 ,
 REGofMAX1DataOut_F3_123, REGofMAX1DataOut_F3_125 , REGofMAX1DataOut_F3_127 , REGofMAX1DataOut_F3_129 , REGofMAX1DataOut_F3_131 , bigaddress222, Super_2_3_2_2_ch3 );
SUPERMUXMODULECONV2_new mux3_1_2_2_ch3 ( REGofMAX1DataOut_F3_37, REGofMAX1DataOut_F3_39 , REGofMAX1DataOut_F3_41 , REGofMAX1DataOut_F3_43 , REGofMAX1DataOut_F3_45 , REGofMAX1DataOut_F3_61 ,
 REGofMAX1DataOut_F3_63 , REGofMAX1DataOut_F3_65 , REGofMAX1DataOut_F3_67 , REGofMAX1DataOut_F3_69 , REGofMAX1DataOut_F3_85 , REGofMAX1DataOut_F3_87 , REGofMAX1DataOut_F3_89 ,
 REGofMAX1DataOut_F3_91, REGofMAX1DataOut_F3_93 , REGofMAX1DataOut_F3_109 , REGofMAX1DataOut_F3_111 , REGofMAX1DataOut_F3_113 , REGofMAX1DataOut_F3_115 , REGofMAX1DataOut_F3_117 ,
 REGofMAX1DataOut_F3_133, REGofMAX1DataOut_F3_135 ,REGofMAX1DataOut_F3_137  , REGofMAX1DataOut_F3_139 , REGofMAX1DataOut_F3_141 , bigaddress222, Super_3_1_2_2_ch3 );
SUPERMUXMODULECONV2_new mux3_2_2_2_ch3 ( REGofMAX1DataOut_F3_38, REGofMAX1DataOut_F3_40 , REGofMAX1DataOut_F3_42 , REGofMAX1DataOut_F3_44 , REGofMAX1DataOut_F3_46 , REGofMAX1DataOut_F3_62 ,
 REGofMAX1DataOut_F3_64 , REGofMAX1DataOut_F3_66 , REGofMAX1DataOut_F3_68 , REGofMAX1DataOut_F3_70 , REGofMAX1DataOut_F3_86 , REGofMAX1DataOut_F3_88 , REGofMAX1DataOut_F3_90 ,
 REGofMAX1DataOut_F3_92, REGofMAX1DataOut_F3_94 , REGofMAX1DataOut_F3_110 , REGofMAX1DataOut_F3_112 , REGofMAX1DataOut_F3_114 , REGofMAX1DataOut_F3_116 , REGofMAX1DataOut_F3_118 ,
REGofMAX1DataOut_F3_134 , REGofMAX1DataOut_F3_136 , REGofMAX1DataOut_F3_138 , REGofMAX1DataOut_F3_140 , REGofMAX1DataOut_F3_142 , bigaddress222, Super_3_2_2_2_ch3 );
SUPERMUXMODULECONV2_new mux3_3_2_2_ch3 ( REGofMAX1DataOut_F3_39, REGofMAX1DataOut_F3_41 , REGofMAX1DataOut_F3_43 , REGofMAX1DataOut_F3_45 , REGofMAX1DataOut_F3_47 , REGofMAX1DataOut_F3_63 ,
 REGofMAX1DataOut_F3_65 , REGofMAX1DataOut_F3_67 , REGofMAX1DataOut_F3_69 , REGofMAX1DataOut_F3_71 , REGofMAX1DataOut_F3_87 , REGofMAX1DataOut_F3_89 , REGofMAX1DataOut_F3_91 ,
 REGofMAX1DataOut_F3_93, REGofMAX1DataOut_F3_95 , REGofMAX1DataOut_F3_111 , REGofMAX1DataOut_F3_113 , REGofMAX1DataOut_F3_115 , REGofMAX1DataOut_F3_117 , REGofMAX1DataOut_F3_119 ,
 REGofMAX1DataOut_F3_135, REGofMAX1DataOut_F3_137 , REGofMAX1DataOut_F3_139 , REGofMAX1DataOut_F3_141 ,  REGofMAX1DataOut_F3_143, bigaddress222, Super_3_3_2_2_ch3 );



MUX9X1_conv2 In3_CONV2_MUX0 ( Super_1_1_1_1_ch3 , Super_1_2_1_1_ch3 , Super_1_3_1_1_ch3 , Super_2_1_1_1_ch3 , Super_2_2_1_1_ch3 , Super_2_3_1_1_ch3 , Super_3_1_1_1_ch3 , Super_3_2_1_1_ch3 , Super_3_3_1_1_ch3  ,  CONV2_address , In3_CONV2_MUXout0 );
MUX9X1_conv2 In3_CONV2_MUX1 ( Super_1_1_1_2_ch3 , Super_1_2_1_2_ch3 , Super_1_3_1_2_ch3 , Super_2_1_1_2_ch3 , Super_2_2_1_2_ch3 , Super_2_3_1_2_ch3 , Super_3_1_1_2_ch3 ,   Super_3_2_1_2_ch3 , Super_3_3_1_2_ch3 ,  CONV2_address , In3_CONV2_MUXout1 );
MUX9X1_conv2 In3_CONV2_MUX10 ( Super_1_1_2_1_ch3 , Super_1_2_2_1_ch3 , Super_1_3_2_1_ch3 , Super_2_1_2_1_ch3 , Super_2_2_2_1_ch3 , Super_2_3_2_1_ch3 , Super_3_1_2_1_ch3 , Super_3_2_2_1_ch3 , Super_3_3_2_1_ch3   ,  CONV2_address , In3_CONV2_MUXout10 );
MUX9X1_conv2 In3_CONV2_MUX11 (  Super_1_1_2_2_ch3 , Super_1_2_2_2_ch3 , Super_1_3_2_2_ch3 , Super_2_1_2_2_ch3 , Super_2_2_2_2_ch3 , Super_2_3_2_2_ch3 , Super_3_1_2_2_ch3 ,  Super_3_2_2_2_ch3 , Super_3_3_2_2_ch3  ,  CONV2_address , In3_CONV2_MUXout11 );



MAC_9 In3_CONV2_MAC0_F1 (In3_CONV2_ROMout, In3_CONV2_MUXout0 , clk, In3_CONV2_MACoutF1_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC1_F1  (In3_CONV2_ROMout, In3_CONV2_MUXout1 , clk, In3_CONV2_MACoutF1_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC10_F1  (In3_CONV2_ROMout, In3_CONV2_MUXout10 , clk, In3_CONV2_MACoutF1_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC11_F1  (In3_CONV2_ROMout, In3_CONV2_MUXout11 , clk, In3_CONV2_MACoutF1_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In3_CONV2_MAC0_F2 (In3_CONV2_ROMout1, In3_CONV2_MUXout0 , clk, In3_CONV2_MACoutF2_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC1_F2  (In3_CONV2_ROMout1, In3_CONV2_MUXout1 , clk, In3_CONV2_MACoutF2_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC10_F2  (In3_CONV2_ROMout1, In3_CONV2_MUXout10 , clk, In3_CONV2_MACoutF2_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC11_F2  (In3_CONV2_ROMout1, In3_CONV2_MUXout11 , clk, In3_CONV2_MACoutF2_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In3_CONV2_MAC0_F3 (In3_CONV2_ROMout2, In3_CONV2_MUXout0 , clk, In3_CONV2_MACoutF3_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC1_F3 (In3_CONV2_ROMout2, In3_CONV2_MUXout1 , clk, In3_CONV2_MACoutF3_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC10_F3 (In3_CONV2_ROMout2, In3_CONV2_MUXout10 , clk, In3_CONV2_MACoutF3_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC11_F3 (In3_CONV2_ROMout2, In3_CONV2_MUXout11 , clk, In3_CONV2_MACoutF3_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In3_CONV2_MAC0_F4 (In3_CONV2_ROMout3, In3_CONV2_MUXout0 , clk, In3_CONV2_MACoutF4_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC1_F4  (In3_CONV2_ROMout3, In3_CONV2_MUXout1 , clk, In3_CONV2_MACoutF4_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC10_F4  (In3_CONV2_ROMout3, In3_CONV2_MUXout10 , clk, In3_CONV2_MACoutF4_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In3_CONV2_MAC11_F4  (In3_CONV2_ROMout3, In3_CONV2_MUXout11 , clk, In3_CONV2_MACoutF4_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);


//input4th channel



SUPERMUXMODULECONV2_new mux1_1_1_1_ch4 ( REGofMAX1DataOut_F4_0, REGofMAX1DataOut_F4_2 , REGofMAX1DataOut_F4_4 , REGofMAX1DataOut_F4_6 , REGofMAX1DataOut_F4_8 , REGofMAX1DataOut_F4_24 ,
 REGofMAX1DataOut_F4_26 , REGofMAX1DataOut_F4_28 , REGofMAX1DataOut_F4_30 , REGofMAX1DataOut_F4_32 , REGofMAX1DataOut_F4_48 , REGofMAX1DataOut_F4_50 , REGofMAX1DataOut_F4_52 ,
 REGofMAX1DataOut_F4_54, REGofMAX1DataOut_F4_56 , REGofMAX1DataOut_F4_72 , REGofMAX1DataOut_F4_74 , REGofMAX1DataOut_F4_76 , REGofMAX1DataOut_F4_78 , REGofMAX1DataOut_F4_80 ,
 REGofMAX1DataOut_F4_96, REGofMAX1DataOut_F4_98 ,REGofMAX1DataOut_F4_100  , REGofMAX1DataOut_F4_102 , REGofMAX1DataOut_F4_104 , bigaddress222, Super_1_1_1_1_ch4 );
SUPERMUXMODULECONV2_new mux1_2_1_1_ch4 ( REGofMAX1DataOut_F4_1 , REGofMAX1DataOut_F4_3 , REGofMAX1DataOut_F4_5 , REGofMAX1DataOut_F4_7 , REGofMAX1DataOut_F4_9 , REGofMAX1DataOut_F4_25 ,
 REGofMAX1DataOut_F4_27 , REGofMAX1DataOut_F4_29 , REGofMAX1DataOut_F4_31 , REGofMAX1DataOut_F4_33 , REGofMAX1DataOut_F4_49 , REGofMAX1DataOut_F4_51 , REGofMAX1DataOut_F4_53 ,
 REGofMAX1DataOut_F4_55, REGofMAX1DataOut_F4_57 , REGofMAX1DataOut_F4_73 , REGofMAX1DataOut_F4_75 , REGofMAX1DataOut_F4_77 , REGofMAX1DataOut_F4_79 , REGofMAX1DataOut_F4_81 ,
 REGofMAX1DataOut_F4_97, REGofMAX1DataOut_F4_99 , REGofMAX1DataOut_F4_101 , REGofMAX1DataOut_F4_103 ,  REGofMAX1DataOut_F4_105, bigaddress222, Super_1_2_1_1_ch4 );
SUPERMUXMODULECONV2_new mux1_3_1_1_ch4 ( REGofMAX1DataOut_F4_2,  REGofMAX1DataOut_F4_4, REGofMAX1DataOut_F4_6 , REGofMAX1DataOut_F4_8 , REGofMAX1DataOut_F4_10 , REGofMAX1DataOut_F4_26 ,
 REGofMAX1DataOut_F4_28 , REGofMAX1DataOut_F4_30 , REGofMAX1DataOut_F4_32 , REGofMAX1DataOut_F4_34 , REGofMAX1DataOut_F4_50 , REGofMAX1DataOut_F4_52 , REGofMAX1DataOut_F4_54 ,
 REGofMAX1DataOut_F4_56, REGofMAX1DataOut_F4_58 , REGofMAX1DataOut_F4_74 , REGofMAX1DataOut_F4_76 , REGofMAX1DataOut_F4_78 , REGofMAX1DataOut_F4_80 , REGofMAX1DataOut_F4_82 ,
 REGofMAX1DataOut_F4_98, REGofMAX1DataOut_F4_100 , REGofMAX1DataOut_F4_102 , REGofMAX1DataOut_F4_104 , REGofMAX1DataOut_F4_106 , bigaddress222, Super_1_3_1_1_ch4 );
SUPERMUXMODULECONV2_new mux2_1_1_1_ch4 ( REGofMAX1DataOut_F4_12 ,REGofMAX1DataOut_F4_14  , REGofMAX1DataOut_F4_16 , REGofMAX1DataOut_F4_18 , REGofMAX1DataOut_F4_20 , REGofMAX1DataOut_F4_36 ,
 REGofMAX1DataOut_F4_38 , REGofMAX1DataOut_F4_40 , REGofMAX1DataOut_F4_42 , REGofMAX1DataOut_F4_44 , REGofMAX1DataOut_F4_60 , REGofMAX1DataOut_F4_62 , REGofMAX1DataOut_F4_64 ,
 REGofMAX1DataOut_F4_66, REGofMAX1DataOut_F4_68 , REGofMAX1DataOut_F4_84 , REGofMAX1DataOut_F4_86 , REGofMAX1DataOut_F4_88 , REGofMAX1DataOut_F4_90 , REGofMAX1DataOut_F4_92  ,
 REGofMAX1DataOut_F4_108, REGofMAX1DataOut_F4_110 , REGofMAX1DataOut_F4_112 , REGofMAX1DataOut_F4_114 , REGofMAX1DataOut_F4_116 , bigaddress222, Super_2_1_1_1_ch4 );
SUPERMUXMODULECONV2_new mux2_2_1_1_ch4 ( REGofMAX1DataOut_F4_13, REGofMAX1DataOut_F4_15 , REGofMAX1DataOut_F4_17 , REGofMAX1DataOut_F4_19 , REGofMAX1DataOut_F4_21 , REGofMAX1DataOut_F4_37 ,
 REGofMAX1DataOut_F4_39 , REGofMAX1DataOut_F4_41 , REGofMAX1DataOut_F4_43 , REGofMAX1DataOut_F4_45 , REGofMAX1DataOut_F4_61 , REGofMAX1DataOut_F4_63 , REGofMAX1DataOut_F4_65 ,
 REGofMAX1DataOut_F4_67, REGofMAX1DataOut_F4_69 , REGofMAX1DataOut_F4_85 , REGofMAX1DataOut_F4_87 , REGofMAX1DataOut_F4_89 , REGofMAX1DataOut_F4_91 ,REGofMAX1DataOut_F4_93  ,
 REGofMAX1DataOut_F4_109, REGofMAX1DataOut_F4_111 , REGofMAX1DataOut_F4_113 , REGofMAX1DataOut_F4_115 ,REGofMAX1DataOut_F4_117  , bigaddress222, Super_2_2_1_1_ch4 );
SUPERMUXMODULECONV2_new mux2_3_1_1_ch4 ( REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_16  , REGofMAX1DataOut_F4_18 , REGofMAX1DataOut_F4_20 , REGofMAX1DataOut_F4_22 , REGofMAX1DataOut_F4_38 ,
 REGofMAX1DataOut_F4_40 , REGofMAX1DataOut_F4_42 , REGofMAX1DataOut_F4_44 , REGofMAX1DataOut_F4_46 , REGofMAX1DataOut_F4_62 , REGofMAX1DataOut_F4_64 , REGofMAX1DataOut_F4_66 ,
 REGofMAX1DataOut_F4_68, REGofMAX1DataOut_F4_70 , REGofMAX1DataOut_F4_86 , REGofMAX1DataOut_F4_88 , REGofMAX1DataOut_F4_90 , REGofMAX1DataOut_F4_92 , REGofMAX1DataOut_F4_94 ,
 REGofMAX1DataOut_F4_110, REGofMAX1DataOut_F4_112 , REGofMAX1DataOut_F4_114 , REGofMAX1DataOut_F4_116 , REGofMAX1DataOut_F4_118 , bigaddress222, Super_2_3_1_1_ch4 );
SUPERMUXMODULECONV2_new mux3_1_1_1_ch4 ( REGofMAX1DataOut_F4_24, REGofMAX1DataOut_F4_26 , REGofMAX1DataOut_F4_28 , REGofMAX1DataOut_F4_30 , REGofMAX1DataOut_F4_32 , REGofMAX1DataOut_F4_48 ,
 REGofMAX1DataOut_F4_50 , REGofMAX1DataOut_F4_52 , REGofMAX1DataOut_F4_54 , REGofMAX1DataOut_F4_56 , REGofMAX1DataOut_F4_72 , REGofMAX1DataOut_F4_74 , REGofMAX1DataOut_F4_76 ,
 REGofMAX1DataOut_F4_78, REGofMAX1DataOut_F4_80 , REGofMAX1DataOut_F4_96 , REGofMAX1DataOut_F4_98 , REGofMAX1DataOut_F4_100 , REGofMAX1DataOut_F4_102 , REGofMAX1DataOut_F4_104 ,
 REGofMAX1DataOut_F4_120, REGofMAX1DataOut_F4_122 , REGofMAX1DataOut_F4_124 , REGofMAX1DataOut_F4_126 , REGofMAX1DataOut_F4_128 , bigaddress222, Super_3_1_1_1_ch4 );
SUPERMUXMODULECONV2_new mux3_2_1_1_ch4 ( REGofMAX1DataOut_F4_25, REGofMAX1DataOut_F4_27 , REGofMAX1DataOut_F4_29 , REGofMAX1DataOut_F4_31 , REGofMAX1DataOut_F4_33 , REGofMAX1DataOut_F4_49 ,
 REGofMAX1DataOut_F4_51 ,REGofMAX1DataOut_F4_53  , REGofMAX1DataOut_F4_55 , REGofMAX1DataOut_F4_57 , REGofMAX1DataOut_F4_73 , REGofMAX1DataOut_F4_75 , REGofMAX1DataOut_F4_77 ,
REGofMAX1DataOut_F4_79 , REGofMAX1DataOut_F4_81 , REGofMAX1DataOut_F4_97 , REGofMAX1DataOut_F4_99 , REGofMAX1DataOut_F4_101 , REGofMAX1DataOut_F4_103 , REGofMAX1DataOut_F4_105 ,
 REGofMAX1DataOut_F4_121 , REGofMAX1DataOut_F4_123 , REGofMAX1DataOut_F4_125 , REGofMAX1DataOut_F4_127 , REGofMAX1DataOut_F4_129 , bigaddress222, Super_3_2_1_1_ch4 );
SUPERMUXMODULECONV2_new mux3_3_1_1_ch4 ( REGofMAX1DataOut_F4_26, REGofMAX1DataOut_F4_28 , REGofMAX1DataOut_F4_30 , REGofMAX1DataOut_F4_32 , REGofMAX1DataOut_F4_34 , REGofMAX1DataOut_F4_50 ,
REGofMAX1DataOut_F4_52  , REGofMAX1DataOut_F4_54 , REGofMAX1DataOut_F4_56 , REGofMAX1DataOut_F4_58 , REGofMAX1DataOut_F4_74 , REGofMAX1DataOut_F4_76 , REGofMAX1DataOut_F4_78 ,
REGofMAX1DataOut_F4_80 , REGofMAX1DataOut_F4_82 , REGofMAX1DataOut_F4_98 , REGofMAX1DataOut_F4_100 , REGofMAX1DataOut_F4_102 , REGofMAX1DataOut_F4_104 , REGofMAX1DataOut_F4_106 ,
 REGofMAX1DataOut_F4_122 , REGofMAX1DataOut_F4_124 , REGofMAX1DataOut_F4_126 , REGofMAX1DataOut_F4_128 , REGofMAX1DataOut_F4_130 , bigaddress222, Super_3_3_1_1_ch4 );



SUPERMUXMODULECONV2_new mux1_1_1_2_ch4 ( REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_3  , REGofMAX1DataOut_F4_5 , REGofMAX1DataOut_F4_7 , REGofMAX1DataOut_F4_9 , REGofMAX1DataOut_F4_25 ,
REGofMAX1DataOut_F4_27 , REGofMAX1DataOut_F4_29 , REGofMAX1DataOut_F4_31 , REGofMAX1DataOut_F4_33 , REGofMAX1DataOut_F4_49 , REGofMAX1DataOut_F4_51 ,REGofMAX1DataOut_F4_53  ,
 REGofMAX1DataOut_F4_55 ,REGofMAX1DataOut_F4_57  , REGofMAX1DataOut_F4_73 , REGofMAX1DataOut_F4_75 , REGofMAX1DataOut_F4_77 , REGofMAX1DataOut_F4_79 , REGofMAX1DataOut_F4_81 ,
 REGofMAX1DataOut_F4_97, REGofMAX1DataOut_F4_99 , REGofMAX1DataOut_F4_101 , REGofMAX1DataOut_F4_103 , REGofMAX1DataOut_F4_105 , bigaddress222, Super_1_1_1_2_ch4 );
SUPERMUXMODULECONV2_new mux1_2_1_2_ch4 ( REGofMAX1DataOut_F4_2, REGofMAX1DataOut_F4_4 , REGofMAX1DataOut_F4_6 , REGofMAX1DataOut_F4_8 , REGofMAX1DataOut_F4_10 , REGofMAX1DataOut_F4_26 ,
REGofMAX1DataOut_F4_28 , REGofMAX1DataOut_F4_30 , REGofMAX1DataOut_F4_32 , REGofMAX1DataOut_F4_34 , REGofMAX1DataOut_F4_50 , REGofMAX1DataOut_F4_52 ,REGofMAX1DataOut_F4_54  ,
 REGofMAX1DataOut_F4_56 , REGofMAX1DataOut_F4_58 , REGofMAX1DataOut_F4_74 , REGofMAX1DataOut_F4_76 , REGofMAX1DataOut_F4_78 , REGofMAX1DataOut_F4_80 , REGofMAX1DataOut_F4_82 ,
 REGofMAX1DataOut_F4_98, REGofMAX1DataOut_F4_100 , REGofMAX1DataOut_F4_102 , REGofMAX1DataOut_F4_104 , REGofMAX1DataOut_F4_106 , bigaddress222, Super_1_2_1_2_ch4 );
SUPERMUXMODULECONV2_new mux1_3_1_2_ch4 ( REGofMAX1DataOut_F4_3, REGofMAX1DataOut_F4_5 , REGofMAX1DataOut_F4_7 , REGofMAX1DataOut_F4_9 , REGofMAX1DataOut_F4_11 , REGofMAX1DataOut_F4_27 ,
REGofMAX1DataOut_F4_29 , REGofMAX1DataOut_F4_31 , REGofMAX1DataOut_F4_33 , REGofMAX1DataOut_F4_35 , REGofMAX1DataOut_F4_51 , REGofMAX1DataOut_F4_53 , REGofMAX1DataOut_F4_55 ,
 REGofMAX1DataOut_F4_57 , REGofMAX1DataOut_F4_59 , REGofMAX1DataOut_F4_75 , REGofMAX1DataOut_F4_77 , REGofMAX1DataOut_F4_79 , REGofMAX1DataOut_F4_81 , REGofMAX1DataOut_F4_83 ,
 REGofMAX1DataOut_F4_99, REGofMAX1DataOut_F4_101 , REGofMAX1DataOut_F4_103 , REGofMAX1DataOut_F4_105 , REGofMAX1DataOut_F4_107 , bigaddress222, Super_1_3_1_2_ch4 );
SUPERMUXMODULECONV2_new mux2_1_1_2_ch4 ( REGofMAX1DataOut_F4_13, REGofMAX1DataOut_F4_15 , REGofMAX1DataOut_F4_17 , REGofMAX1DataOut_F4_19 , REGofMAX1DataOut_F4_21 , REGofMAX1DataOut_F4_37 ,
REGofMAX1DataOut_F4_39 , REGofMAX1DataOut_F4_41 , REGofMAX1DataOut_F4_43 , REGofMAX1DataOut_F4_45 , REGofMAX1DataOut_F4_61 , REGofMAX1DataOut_F4_63  ,REGofMAX1DataOut_F4_65  ,
 REGofMAX1DataOut_F4_67 , REGofMAX1DataOut_F4_69 , REGofMAX1DataOut_F4_85 , REGofMAX1DataOut_F4_87 , REGofMAX1DataOut_F4_89 , REGofMAX1DataOut_F4_91 , REGofMAX1DataOut_F4_93 ,
 REGofMAX1DataOut_F4_109, REGofMAX1DataOut_F4_111 , REGofMAX1DataOut_F4_113 , REGofMAX1DataOut_F4_115 , REGofMAX1DataOut_F4_117 , bigaddress222, Super_2_1_1_2_ch4 );
SUPERMUXMODULECONV2_new mux2_2_1_2_ch4 ( REGofMAX1DataOut_F4_14, REGofMAX1DataOut_F4_16 , REGofMAX1DataOut_F4_18 , REGofMAX1DataOut_F4_20 , REGofMAX1DataOut_F4_22 , REGofMAX1DataOut_F4_38 ,
REGofMAX1DataOut_F4_40  , REGofMAX1DataOut_F4_42 , REGofMAX1DataOut_F4_44 , REGofMAX1DataOut_F4_46 , REGofMAX1DataOut_F4_62 , REGofMAX1DataOut_F4_64 ,REGofMAX1DataOut_F4_66  ,
 REGofMAX1DataOut_F4_68 , REGofMAX1DataOut_F4_70 , REGofMAX1DataOut_F4_86 , REGofMAX1DataOut_F4_88 , REGofMAX1DataOut_F4_90 , REGofMAX1DataOut_F4_92 , REGofMAX1DataOut_F4_94 ,
 REGofMAX1DataOut_F4_110, REGofMAX1DataOut_F4_112 , REGofMAX1DataOut_F4_114 , REGofMAX1DataOut_F4_116 , REGofMAX1DataOut_F4_118 , bigaddress222, Super_2_2_1_2_ch4 );
SUPERMUXMODULECONV2_new mux2_3_1_2_ch4 ( REGofMAX1DataOut_F4_15, REGofMAX1DataOut_F4_17 , REGofMAX1DataOut_F4_19 , REGofMAX1DataOut_F4_21 , REGofMAX1DataOut_F4_23 , REGofMAX1DataOut_F4_39 ,
REGofMAX1DataOut_F4_41  , REGofMAX1DataOut_F4_43 , REGofMAX1DataOut_F4_45 , REGofMAX1DataOut_F4_47 , REGofMAX1DataOut_F4_63 , REGofMAX1DataOut_F4_65 ,REGofMAX1DataOut_F4_67  ,
 REGofMAX1DataOut_F4_69 , REGofMAX1DataOut_F4_71 , REGofMAX1DataOut_F4_87 , REGofMAX1DataOut_F4_89 , REGofMAX1DataOut_F4_91 , REGofMAX1DataOut_F4_93 , REGofMAX1DataOut_F4_95 ,
 REGofMAX1DataOut_F4_111, REGofMAX1DataOut_F4_113 , REGofMAX1DataOut_F4_115 , REGofMAX1DataOut_F4_117 , REGofMAX1DataOut_F4_119 , bigaddress222, Super_2_3_1_2_ch4 );
SUPERMUXMODULECONV2_new mux3_1_1_2_ch4 ( REGofMAX1DataOut_F4_25, REGofMAX1DataOut_F4_27 , REGofMAX1DataOut_F4_29 , REGofMAX1DataOut_F4_31 , REGofMAX1DataOut_F4_33 , REGofMAX1DataOut_F4_49 ,
REGofMAX1DataOut_F4_51 , REGofMAX1DataOut_F4_53 , REGofMAX1DataOut_F4_55 , REGofMAX1DataOut_F4_57 , REGofMAX1DataOut_F4_73 , REGofMAX1DataOut_F4_75 ,REGofMAX1DataOut_F4_77  ,
 REGofMAX1DataOut_F4_79 , REGofMAX1DataOut_F4_81 , REGofMAX1DataOut_F4_97 , REGofMAX1DataOut_F4_99 , REGofMAX1DataOut_F4_101 , REGofMAX1DataOut_F4_103 , REGofMAX1DataOut_F4_105 ,
REGofMAX1DataOut_F4_121 , REGofMAX1DataOut_F4_123 , REGofMAX1DataOut_F4_125 , REGofMAX1DataOut_F4_127 , REGofMAX1DataOut_F4_129 , bigaddress222, Super_3_1_1_2_ch4 );
SUPERMUXMODULECONV2_new mux3_2_1_2_ch4 ( REGofMAX1DataOut_F4_26, REGofMAX1DataOut_F4_28 , REGofMAX1DataOut_F4_30 , REGofMAX1DataOut_F4_32 , REGofMAX1DataOut_F4_34 , REGofMAX1DataOut_F4_50 ,
REGofMAX1DataOut_F4_52  , REGofMAX1DataOut_F4_54 , REGofMAX1DataOut_F4_56 , REGofMAX1DataOut_F4_58 , REGofMAX1DataOut_F4_74 , REGofMAX1DataOut_F4_76 ,REGofMAX1DataOut_F4_78  ,
 REGofMAX1DataOut_F4_80 , REGofMAX1DataOut_F4_82 , REGofMAX1DataOut_F4_98 , REGofMAX1DataOut_F4_100 , REGofMAX1DataOut_F4_102 , REGofMAX1DataOut_F4_104 ,REGofMAX1DataOut_F4_106  ,
 REGofMAX1DataOut_F4_122, REGofMAX1DataOut_F4_124 , REGofMAX1DataOut_F4_126 , REGofMAX1DataOut_F4_128 , REGofMAX1DataOut_F4_130 , bigaddress222, Super_3_2_1_2_ch4 );
SUPERMUXMODULECONV2_new mux3_3_1_2_ch4 ( REGofMAX1DataOut_F4_27, REGofMAX1DataOut_F4_29 , REGofMAX1DataOut_F4_31 , REGofMAX1DataOut_F4_33 , REGofMAX1DataOut_F4_35 , REGofMAX1DataOut_F4_51 ,
REGofMAX1DataOut_F4_53 , REGofMAX1DataOut_F4_55 , REGofMAX1DataOut_F4_57 , REGofMAX1DataOut_F4_59 , REGofMAX1DataOut_F4_75 , REGofMAX1DataOut_F4_77 , REGofMAX1DataOut_F4_79 ,
 REGofMAX1DataOut_F4_81 , REGofMAX1DataOut_F4_83 ,REGofMAX1DataOut_F4_99  , REGofMAX1DataOut_F4_101 , REGofMAX1DataOut_F4_103 , REGofMAX1DataOut_F4_105 , REGofMAX1DataOut_F4_107 ,
 REGofMAX1DataOut_F4_123, REGofMAX1DataOut_F4_125 , REGofMAX1DataOut_F4_127 , REGofMAX1DataOut_F4_129 , REGofMAX1DataOut_F4_131 , bigaddress222, Super_3_3_1_2_ch4 );


SUPERMUXMODULECONV2_new mux1_1_2_1_ch4 ( REGofMAX1DataOut_F4_12, REGofMAX1DataOut_F4_14 , REGofMAX1DataOut_F4_16 , REGofMAX1DataOut_F4_18 , REGofMAX1DataOut_F4_20 , REGofMAX1DataOut_F4_36 ,
 REGofMAX1DataOut_F4_38 , REGofMAX1DataOut_F4_40 , REGofMAX1DataOut_F4_42 , REGofMAX1DataOut_F4_44 , REGofMAX1DataOut_F4_60 , REGofMAX1DataOut_F4_62 , REGofMAX1DataOut_F4_64 ,
 REGofMAX1DataOut_F4_66, REGofMAX1DataOut_F4_68 , REGofMAX1DataOut_F4_84 , REGofMAX1DataOut_F4_86 , REGofMAX1DataOut_F4_88 , REGofMAX1DataOut_F4_90 , REGofMAX1DataOut_F4_92 ,
 REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_110  , REGofMAX1DataOut_F4_112 , REGofMAX1DataOut_F4_114 , REGofMAX1DataOut_F4_116 , bigaddress222, Super_1_1_2_1_ch4 );
SUPERMUXMODULECONV2_new mux1_2_2_1_ch4 ( REGofMAX1DataOut_F4_13, REGofMAX1DataOut_F4_15 , REGofMAX1DataOut_F4_17 , REGofMAX1DataOut_F4_19 , REGofMAX1DataOut_F4_21 , REGofMAX1DataOut_F4_37 ,
 REGofMAX1DataOut_F4_39 , REGofMAX1DataOut_F4_41 , REGofMAX1DataOut_F4_43 , REGofMAX1DataOut_F4_45 , REGofMAX1DataOut_F4_61 , REGofMAX1DataOut_F4_63 , REGofMAX1DataOut_F4_65 ,
 REGofMAX1DataOut_F4_67, REGofMAX1DataOut_F4_69 , REGofMAX1DataOut_F4_85 , REGofMAX1DataOut_F4_87 , REGofMAX1DataOut_F4_89 , REGofMAX1DataOut_F4_91 , REGofMAX1DataOut_F4_93 ,
 REGofMAX1DataOut_F4_109, REGofMAX1DataOut_F4_111 , REGofMAX1DataOut_F4_113 , REGofMAX1DataOut_F4_115 , REGofMAX1DataOut_F4_117 , bigaddress222, Super_1_2_2_1_ch4 );
SUPERMUXMODULECONV2_new mux1_3_2_1_ch4 ( REGofMAX1DataOut_F4_14, REGofMAX1DataOut_F4_16 , REGofMAX1DataOut_F4_18 , REGofMAX1DataOut_F4_20 , REGofMAX1DataOut_F4_22 , REGofMAX1DataOut_F4_38 ,
REGofMAX1DataOut_F4_40  , REGofMAX1DataOut_F4_42 , REGofMAX1DataOut_F4_44 , REGofMAX1DataOut_F4_46 , REGofMAX1DataOut_F4_62 , REGofMAX1DataOut_F4_64 ,REGofMAX1DataOut_F4_66 ,
 REGofMAX1DataOut_F4_68 , REGofMAX1DataOut_F4_70 , REGofMAX1DataOut_F4_86 , REGofMAX1DataOut_F4_88 ,REGofMAX1DataOut_F4_90  , REGofMAX1DataOut_F4_92 , REGofMAX1DataOut_F4_94 ,
REGofMAX1DataOut_F4_110 , REGofMAX1DataOut_F4_112 , REGofMAX1DataOut_F4_114 , REGofMAX1DataOut_F4_116 , REGofMAX1DataOut_F4_118 , bigaddress222, Super_1_3_2_1_ch4 );
SUPERMUXMODULECONV2_new mux2_1_2_1_ch4 ( REGofMAX1DataOut_F4_24, REGofMAX1DataOut_F4_26 , REGofMAX1DataOut_F4_28 , REGofMAX1DataOut_F4_30 , REGofMAX1DataOut_F4_32 , REGofMAX1DataOut_F4_48 ,
 REGofMAX1DataOut_F4_50 , REGofMAX1DataOut_F4_52 , REGofMAX1DataOut_F4_54 , REGofMAX1DataOut_F4_56 , REGofMAX1DataOut_F4_72 , REGofMAX1DataOut_F4_74 ,REGofMAX1DataOut_F4_76  ,
 REGofMAX1DataOut_F4_78, REGofMAX1DataOut_F4_80 , REGofMAX1DataOut_F4_96 , REGofMAX1DataOut_F4_98 , REGofMAX1DataOut_F4_100 , REGofMAX1DataOut_F4_102 , REGofMAX1DataOut_F4_104 ,
REGofMAX1DataOut_F4_120 , REGofMAX1DataOut_F4_122 , REGofMAX1DataOut_F4_124 , REGofMAX1DataOut_F4_126 , REGofMAX1DataOut_F4_128 , bigaddress222, Super_2_1_2_1_ch4 );
SUPERMUXMODULECONV2_new mux2_2_2_1_ch4 ( REGofMAX1DataOut_F4_25, REGofMAX1DataOut_F4_27 , REGofMAX1DataOut_F4_29 , REGofMAX1DataOut_F4_31 , REGofMAX1DataOut_F4_33 , REGofMAX1DataOut_F4_49 ,
 REGofMAX1DataOut_F4_51 , REGofMAX1DataOut_F4_53 , REGofMAX1DataOut_F4_55 , REGofMAX1DataOut_F4_57 , REGofMAX1DataOut_F4_73 , REGofMAX1DataOut_F4_75 , REGofMAX1DataOut_F4_77 ,
 REGofMAX1DataOut_F4_79, REGofMAX1DataOut_F4_81 , REGofMAX1DataOut_F4_97 , REGofMAX1DataOut_F4_99 , REGofMAX1DataOut_F4_101 , REGofMAX1DataOut_F4_103 , REGofMAX1DataOut_F4_105 ,
REGofMAX1DataOut_F4_121 , REGofMAX1DataOut_F4_123 , REGofMAX1DataOut_F4_125 , REGofMAX1DataOut_F4_127 , REGofMAX1DataOut_F4_129 , bigaddress222, Super_2_2_2_1_ch4 );
SUPERMUXMODULECONV2_new mux2_3_2_1_ch4 ( REGofMAX1DataOut_F4_26, REGofMAX1DataOut_F4_28 , REGofMAX1DataOut_F4_30 , REGofMAX1DataOut_F4_32 , REGofMAX1DataOut_F4_34 , REGofMAX1DataOut_F4_50 ,
 REGofMAX1DataOut_F4_52 , REGofMAX1DataOut_F4_54 , REGofMAX1DataOut_F4_56 , REGofMAX1DataOut_F4_58 , REGofMAX1DataOut_F4_74 , REGofMAX1DataOut_F4_76 ,REGofMAX1DataOut_F4_78  ,
 REGofMAX1DataOut_F4_80, REGofMAX1DataOut_F4_82 , REGofMAX1DataOut_F4_98 , REGofMAX1DataOut_F4_100 , REGofMAX1DataOut_F4_102 , REGofMAX1DataOut_F4_104 , REGofMAX1DataOut_F4_106 ,
 REGofMAX1DataOut_F4_122, REGofMAX1DataOut_F4_124 , REGofMAX1DataOut_F4_126 , REGofMAX1DataOut_F4_128 , REGofMAX1DataOut_F4_130 , bigaddress222, Super_2_3_2_1_ch4 );
SUPERMUXMODULECONV2_new mux3_1_2_1_ch4 ( REGofMAX1DataOut_F4_36, REGofMAX1DataOut_F4_38 , REGofMAX1DataOut_F4_40 , REGofMAX1DataOut_F4_42 , REGofMAX1DataOut_F4_44 , REGofMAX1DataOut_F4_60 ,
 REGofMAX1DataOut_F4_62 , REGofMAX1DataOut_F4_64 , REGofMAX1DataOut_F4_66 , REGofMAX1DataOut_F4_68 , REGofMAX1DataOut_F4_84 , REGofMAX1DataOut_F4_86 ,REGofMAX1DataOut_F4_88  ,
 REGofMAX1DataOut_F4_90, REGofMAX1DataOut_F4_92 , REGofMAX1DataOut_F4_108 , REGofMAX1DataOut_F4_110 , REGofMAX1DataOut_F4_112 , REGofMAX1DataOut_F4_114 , REGofMAX1DataOut_F4_116 ,
 REGofMAX1DataOut_F4_132, REGofMAX1DataOut_F4_134 , REGofMAX1DataOut_F4_136 , REGofMAX1DataOut_F4_138 , REGofMAX1DataOut_F4_140 , bigaddress222, Super_3_1_2_1_ch4 );
SUPERMUXMODULECONV2_new mux3_2_2_1_ch4 ( REGofMAX1DataOut_F4_37, REGofMAX1DataOut_F4_39 , REGofMAX1DataOut_F4_41 , REGofMAX1DataOut_F4_43 , REGofMAX1DataOut_F4_45 , REGofMAX1DataOut_F4_61 ,
 REGofMAX1DataOut_F4_63 , REGofMAX1DataOut_F4_65 , REGofMAX1DataOut_F4_67 , REGofMAX1DataOut_F4_69 , REGofMAX1DataOut_F4_85 , REGofMAX1DataOut_F4_87 , REGofMAX1DataOut_F4_89 ,
 REGofMAX1DataOut_F4_91, REGofMAX1DataOut_F4_93 , REGofMAX1DataOut_F4_109 , REGofMAX1DataOut_F4_111 , REGofMAX1DataOut_F4_113 , REGofMAX1DataOut_F4_115 , REGofMAX1DataOut_F4_117 ,
 REGofMAX1DataOut_F4_133, REGofMAX1DataOut_F4_135 , REGofMAX1DataOut_F4_137 , REGofMAX1DataOut_F4_139 , REGofMAX1DataOut_F4_141 , bigaddress222, Super_3_2_2_1_ch4 );
SUPERMUXMODULECONV2_new mux3_3_2_1_ch4 ( REGofMAX1DataOut_F4_38, REGofMAX1DataOut_F4_40 , REGofMAX1DataOut_F4_42 , REGofMAX1DataOut_F4_44 , REGofMAX1DataOut_F4_46 , REGofMAX1DataOut_F4_62 ,
 REGofMAX1DataOut_F4_64 , REGofMAX1DataOut_F4_66 , REGofMAX1DataOut_F4_68 , REGofMAX1DataOut_F4_70 , REGofMAX1DataOut_F4_86 , REGofMAX1DataOut_F4_88 , REGofMAX1DataOut_F4_90 ,
 REGofMAX1DataOut_F4_92, REGofMAX1DataOut_F4_94 , REGofMAX1DataOut_F4_110 , REGofMAX1DataOut_F4_112 , REGofMAX1DataOut_F4_114 , REGofMAX1DataOut_F4_116 , REGofMAX1DataOut_F4_118 ,
 REGofMAX1DataOut_F4_134,  REGofMAX1DataOut_F4_136, REGofMAX1DataOut_F4_138 , REGofMAX1DataOut_F4_140 , REGofMAX1DataOut_F4_142 , bigaddress222, Super_3_3_2_1_ch4 );


SUPERMUXMODULECONV2_new mux1_1_2_2_ch4 ( REGofMAX1DataOut_F4_13, REGofMAX1DataOut_F4_15 , REGofMAX1DataOut_F4_17 , REGofMAX1DataOut_F4_19 , REGofMAX1DataOut_F4_21 , REGofMAX1DataOut_F4_37 ,
 REGofMAX1DataOut_F4_39 , REGofMAX1DataOut_F4_41 , REGofMAX1DataOut_F4_43 , REGofMAX1DataOut_F4_45 , REGofMAX1DataOut_F4_61 , REGofMAX1DataOut_F4_63 , REGofMAX1DataOut_F4_65 ,
 REGofMAX1DataOut_F4_67, REGofMAX1DataOut_F4_69 , REGofMAX1DataOut_F4_85 , REGofMAX1DataOut_F4_87 , REGofMAX1DataOut_F4_89 , REGofMAX1DataOut_F4_91 , REGofMAX1DataOut_F4_93 ,
 REGofMAX1DataOut_F4_109, REGofMAX1DataOut_F4_111 , REGofMAX1DataOut_F4_113 , REGofMAX1DataOut_F4_115 , REGofMAX1DataOut_F4_117 , bigaddress222, Super_1_1_2_2_ch4 );
SUPERMUXMODULECONV2_new mux1_2_2_2_ch4 ( REGofMAX1DataOut_F4_14, REGofMAX1DataOut_F4_16 , REGofMAX1DataOut_F4_18 , REGofMAX1DataOut_F4_20 , REGofMAX1DataOut_F4_22 , REGofMAX1DataOut_F4_38 ,
 REGofMAX1DataOut_F4_40 , REGofMAX1DataOut_F4_42 , REGofMAX1DataOut_F4_44 , REGofMAX1DataOut_F4_46 , REGofMAX1DataOut_F4_62 , REGofMAX1DataOut_F4_64 , REGofMAX1DataOut_F4_66 ,
REGofMAX1DataOut_F4_68 , REGofMAX1DataOut_F4_70 , REGofMAX1DataOut_F4_86 , REGofMAX1DataOut_F4_88 , REGofMAX1DataOut_F4_90 , REGofMAX1DataOut_F4_92 , REGofMAX1DataOut_F4_94 ,
 REGofMAX1DataOut_F4_110 , REGofMAX1DataOut_F4_112 , REGofMAX1DataOut_F4_114 , REGofMAX1DataOut_F4_116 , REGofMAX1DataOut_F4_118 , bigaddress222, Super_1_2_2_2_ch4 );
SUPERMUXMODULECONV2_new mux1_3_2_2_ch4 ( REGofMAX1DataOut_F4_15, REGofMAX1DataOut_F4_17 , REGofMAX1DataOut_F4_19 , REGofMAX1DataOut_F4_21 , REGofMAX1DataOut_F4_23 , REGofMAX1DataOut_F4_39 ,
 REGofMAX1DataOut_F4_41 , REGofMAX1DataOut_F4_43 , REGofMAX1DataOut_F4_45 , REGofMAX1DataOut_F4_47 , REGofMAX1DataOut_F4_63 , REGofMAX1DataOut_F4_65 , REGofMAX1DataOut_F4_67 ,
 REGofMAX1DataOut_F4_69, REGofMAX1DataOut_F4_71 , REGofMAX1DataOut_F4_87 , REGofMAX1DataOut_F4_89 , REGofMAX1DataOut_F4_91 , REGofMAX1DataOut_F4_93 , REGofMAX1DataOut_F4_95 ,
 REGofMAX1DataOut_F4_111, REGofMAX1DataOut_F4_113 , REGofMAX1DataOut_F4_115 , REGofMAX1DataOut_F4_117 , REGofMAX1DataOut_F4_119 , bigaddress222, Super_1_3_2_2_ch4 );
SUPERMUXMODULECONV2_new mux2_1_2_2_ch4 ( REGofMAX1DataOut_F4_25, REGofMAX1DataOut_F4_27 , REGofMAX1DataOut_F4_29 , REGofMAX1DataOut_F4_31 , REGofMAX1DataOut_F4_33 , REGofMAX1DataOut_F4_49 ,
 REGofMAX1DataOut_F4_51 , REGofMAX1DataOut_F4_53 , REGofMAX1DataOut_F4_55 , REGofMAX1DataOut_F4_57 , REGofMAX1DataOut_F4_73 , REGofMAX1DataOut_F4_75 , REGofMAX1DataOut_F4_77 ,
 REGofMAX1DataOut_F4_79, REGofMAX1DataOut_F4_81 , REGofMAX1DataOut_F4_97 , REGofMAX1DataOut_F4_99 , REGofMAX1DataOut_F4_101 , REGofMAX1DataOut_F4_103 , REGofMAX1DataOut_F4_105 ,
 REGofMAX1DataOut_F4_121, REGofMAX1DataOut_F4_123 , REGofMAX1DataOut_F4_125 , REGofMAX1DataOut_F4_127 , REGofMAX1DataOut_F4_129 , bigaddress222, Super_2_1_2_2_ch4 );
SUPERMUXMODULECONV2_new mux2_2_2_2_ch4 ( REGofMAX1DataOut_F4_26, REGofMAX1DataOut_F4_28 , REGofMAX1DataOut_F4_30 , REGofMAX1DataOut_F4_32 , REGofMAX1DataOut_F4_34 , REGofMAX1DataOut_F4_50 ,
 REGofMAX1DataOut_F4_52 , REGofMAX1DataOut_F4_54 , REGofMAX1DataOut_F4_56 , REGofMAX1DataOut_F4_58 , REGofMAX1DataOut_F4_74 , REGofMAX1DataOut_F4_76 , REGofMAX1DataOut_F4_78 ,
 REGofMAX1DataOut_F4_80, REGofMAX1DataOut_F4_82 , REGofMAX1DataOut_F4_98 , REGofMAX1DataOut_F4_100 , REGofMAX1DataOut_F4_102 , REGofMAX1DataOut_F4_104 , REGofMAX1DataOut_F4_106 ,
 REGofMAX1DataOut_F4_122, REGofMAX1DataOut_F4_124 , REGofMAX1DataOut_F4_126 , REGofMAX1DataOut_F4_128 , REGofMAX1DataOut_F4_130 , bigaddress222, Super_2_2_2_2_ch4 );
SUPERMUXMODULECONV2_new mux2_3_2_2_ch4 ( REGofMAX1DataOut_F4_27, REGofMAX1DataOut_F4_29 , REGofMAX1DataOut_F4_31 , REGofMAX1DataOut_F4_33 , REGofMAX1DataOut_F4_35 , REGofMAX1DataOut_F4_51 ,
 REGofMAX1DataOut_F4_53 , REGofMAX1DataOut_F4_55 , REGofMAX1DataOut_F4_57 , REGofMAX1DataOut_F4_59 , REGofMAX1DataOut_F4_75 , REGofMAX1DataOut_F4_77 , REGofMAX1DataOut_F4_79 ,
 REGofMAX1DataOut_F4_81, REGofMAX1DataOut_F4_83 , REGofMAX1DataOut_F4_99 , REGofMAX1DataOut_F4_101 , REGofMAX1DataOut_F4_103 , REGofMAX1DataOut_F4_105 , REGofMAX1DataOut_F4_107 ,
 REGofMAX1DataOut_F4_123, REGofMAX1DataOut_F4_125 , REGofMAX1DataOut_F4_127 , REGofMAX1DataOut_F4_129 , REGofMAX1DataOut_F4_131 , bigaddress222, Super_2_3_2_2_ch4 );
SUPERMUXMODULECONV2_new mux3_1_2_2_ch4 ( REGofMAX1DataOut_F4_37, REGofMAX1DataOut_F4_39 , REGofMAX1DataOut_F4_41 , REGofMAX1DataOut_F4_43 , REGofMAX1DataOut_F4_45 , REGofMAX1DataOut_F4_61 ,
 REGofMAX1DataOut_F4_63 , REGofMAX1DataOut_F4_65 , REGofMAX1DataOut_F4_67 , REGofMAX1DataOut_F4_69 , REGofMAX1DataOut_F4_85 , REGofMAX1DataOut_F4_87 , REGofMAX1DataOut_F4_89 ,
 REGofMAX1DataOut_F4_91, REGofMAX1DataOut_F4_93 , REGofMAX1DataOut_F4_109 , REGofMAX1DataOut_F4_111 , REGofMAX1DataOut_F4_113 , REGofMAX1DataOut_F4_115 , REGofMAX1DataOut_F4_117 ,
 REGofMAX1DataOut_F4_133, REGofMAX1DataOut_F4_135 ,REGofMAX1DataOut_F4_137  , REGofMAX1DataOut_F4_139 , REGofMAX1DataOut_F4_141 , bigaddress222, Super_3_1_2_2_ch4 );
SUPERMUXMODULECONV2_new mux3_2_2_2_ch4 ( REGofMAX1DataOut_F4_38, REGofMAX1DataOut_F4_40 , REGofMAX1DataOut_F4_42 , REGofMAX1DataOut_F4_44 , REGofMAX1DataOut_F4_46 , REGofMAX1DataOut_F4_62 ,
 REGofMAX1DataOut_F4_64 , REGofMAX1DataOut_F4_66 , REGofMAX1DataOut_F4_68 , REGofMAX1DataOut_F4_70 , REGofMAX1DataOut_F4_86 , REGofMAX1DataOut_F4_88 , REGofMAX1DataOut_F4_90 ,
 REGofMAX1DataOut_F4_92, REGofMAX1DataOut_F4_94 , REGofMAX1DataOut_F4_110 , REGofMAX1DataOut_F4_112 , REGofMAX1DataOut_F4_114 , REGofMAX1DataOut_F4_116 , REGofMAX1DataOut_F4_118 ,
REGofMAX1DataOut_F4_134 , REGofMAX1DataOut_F4_136 , REGofMAX1DataOut_F4_138 , REGofMAX1DataOut_F4_140 , REGofMAX1DataOut_F4_142 , bigaddress222, Super_3_2_2_2_ch4 );
SUPERMUXMODULECONV2_new mux3_3_2_2_ch4 ( REGofMAX1DataOut_F4_39, REGofMAX1DataOut_F4_41 , REGofMAX1DataOut_F4_43 , REGofMAX1DataOut_F4_45 , REGofMAX1DataOut_F4_47 , REGofMAX1DataOut_F4_63 ,
 REGofMAX1DataOut_F4_65 , REGofMAX1DataOut_F4_67 , REGofMAX1DataOut_F4_69 , REGofMAX1DataOut_F4_71 , REGofMAX1DataOut_F4_87 , REGofMAX1DataOut_F4_89 , REGofMAX1DataOut_F4_91 ,
 REGofMAX1DataOut_F4_93, REGofMAX1DataOut_F4_95 , REGofMAX1DataOut_F4_111 , REGofMAX1DataOut_F4_113 , REGofMAX1DataOut_F4_115 , REGofMAX1DataOut_F4_117 , REGofMAX1DataOut_F4_119 ,
 REGofMAX1DataOut_F4_135, REGofMAX1DataOut_F4_137 , REGofMAX1DataOut_F4_139 , REGofMAX1DataOut_F4_141 ,  REGofMAX1DataOut_F4_143, bigaddress222, Super_3_3_2_2_ch4 );



MUX9X1_conv2 In4_CONV2_MUX0 ( Super_1_1_1_1_ch4 , Super_1_2_1_1_ch4 , Super_1_3_1_1_ch4 , Super_2_1_1_1_ch4 , Super_2_2_1_1_ch4 , Super_2_3_1_1_ch4 , Super_3_1_1_1_ch4 , Super_3_2_1_1_ch4 , Super_3_3_1_1_ch4  ,  CONV2_address , In4_CONV2_MUXout0 );
MUX9X1_conv2 In4_CONV2_MUX1 ( Super_1_1_1_2_ch4 , Super_1_2_1_2_ch4 , Super_1_3_1_2_ch4 , Super_2_1_1_2_ch4 , Super_2_2_1_2_ch4 , Super_2_3_1_2_ch4 , Super_3_1_1_2_ch4 ,   Super_3_2_1_2_ch4 , Super_3_3_1_2_ch4 ,  CONV2_address , In4_CONV2_MUXout1 );
MUX9X1_conv2 In4_CONV2_MUX10 ( Super_1_1_2_1_ch4 , Super_1_2_2_1_ch4 , Super_1_3_2_1_ch4 , Super_2_1_2_1_ch4 , Super_2_2_2_1_ch4 , Super_2_3_2_1_ch4 , Super_3_1_2_1_ch4 , Super_3_2_2_1_ch4 , Super_3_3_2_1_ch4   ,  CONV2_address , In4_CONV2_MUXout10 );
MUX9X1_conv2 In4_CONV2_MUX11 (  Super_1_1_2_2_ch4 , Super_1_2_2_2_ch4 , Super_1_3_2_2_ch4 , Super_2_1_2_2_ch4 , Super_2_2_2_2_ch4 , Super_2_3_2_2_ch4 , Super_3_1_2_2_ch4 ,  Super_3_2_2_2_ch4 , Super_3_3_2_2_ch4  ,  CONV2_address , In4_CONV2_MUXout11 );



MAC_9 In4_CONV2_MAC0_F1 (In4_CONV2_ROMout, In4_CONV2_MUXout0 , clk, In4_CONV2_MACoutF1_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC1_F1  (In4_CONV2_ROMout, In4_CONV2_MUXout1 , clk, In4_CONV2_MACoutF1_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC10_F1  (In4_CONV2_ROMout, In4_CONV2_MUXout10 , clk, In4_CONV2_MACoutF1_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC11_F1  (In4_CONV2_ROMout, In4_CONV2_MUXout11 , clk, In4_CONV2_MACoutF1_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In4_CONV2_MAC0_F2 (In4_CONV2_ROMout1, In4_CONV2_MUXout0 , clk, In4_CONV2_MACoutF2_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC1_F2  (In4_CONV2_ROMout1, In4_CONV2_MUXout1 , clk, In4_CONV2_MACoutF2_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC10_F2  (In4_CONV2_ROMout1, In4_CONV2_MUXout10 , clk, In4_CONV2_MACoutF2_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC11_F2  (In4_CONV2_ROMout1, In4_CONV2_MUXout11 , clk, In4_CONV2_MACoutF2_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In4_CONV2_MAC0_F3 (In4_CONV2_ROMout2, In4_CONV2_MUXout0 , clk, In4_CONV2_MACoutF3_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC1_F3 (In4_CONV2_ROMout2, In4_CONV2_MUXout1 , clk, In4_CONV2_MACoutF3_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC10_F3 (In4_CONV2_ROMout2, In4_CONV2_MUXout10 , clk, In4_CONV2_MACoutF3_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC11_F3 (In4_CONV2_ROMout2, In4_CONV2_MUXout11 , clk, In4_CONV2_MACoutF3_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);

MAC_9 In4_CONV2_MAC0_F4 (In4_CONV2_ROMout3, In4_CONV2_MUXout0 , clk, In4_CONV2_MACoutF4_0 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC1_F4  (In4_CONV2_ROMout3, In4_CONV2_MUXout1 , clk, In4_CONV2_MACoutF4_1 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC10_F4  (In4_CONV2_ROMout3, In4_CONV2_MUXout10 , clk, In4_CONV2_MACoutF4_10 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);
MAC_9 In4_CONV2_MAC11_F4  (In4_CONV2_ROMout3, In4_CONV2_MUXout11 , clk, In4_CONV2_MACoutF4_11 , CONV2_MAC_start, CONV2_MAC_end, resetTheCounter);


wire [6:0] count_3bits; //no ok
wire RST65;
assign  RST65=  (CONV2_counter == 157) ?1'b1 :1'b0; //157
COUNTER_LAYER_65_cycles secondStageCONV2_counter (clk,RST65, count_3bits, LayerStartStage2,tttt);

wire [65:0] CONV2_Final_CONV2_MUXout_F1_0,CONV2_Final_CONV2_MUXout_F1_1,CONV2_Final_CONV2_MUXout_F1_10,CONV2_Final_CONV2_MUXout_F1_11;
wire [65:0] CONV2_Final_CONV2_MUXout_F2_0,CONV2_Final_CONV2_MUXout_F2_1,CONV2_Final_CONV2_MUXout_F2_10,CONV2_Final_CONV2_MUXout_F2_11;
wire [65:0] CONV2_Final_CONV2_MUXout_F3_0,CONV2_Final_CONV2_MUXout_F3_1,CONV2_Final_CONV2_MUXout_F3_10,CONV2_Final_CONV2_MUXout_F3_11;
wire [65:0] CONV2_Final_CONV2_MUXout_F4_0,CONV2_Final_CONV2_MUXout_F4_1,CONV2_Final_CONV2_MUXout_F4_10,CONV2_Final_CONV2_MUXout_F4_11;



MUX5X1_13 F1_0 (In1_CONV2_MACoutF1_0  , In2_CONV2_MACoutF1_0  , In3_CONV2_MACoutF1_0  , In4_CONV2_MACoutF1_0  , Filter1BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F1_0 );
MUX5X1_13 F1_1 (In1_CONV2_MACoutF1_1  , In2_CONV2_MACoutF1_1  , In3_CONV2_MACoutF1_1  , In4_CONV2_MACoutF1_1  , Filter1BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F1_1 );
MUX5X1_13 F1_10 (In1_CONV2_MACoutF1_10  , In2_CONV2_MACoutF1_10  , In3_CONV2_MACoutF1_10  , In4_CONV2_MACoutF1_10  , Filter1BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F1_10 );
MUX5X1_13 F1_11 (In1_CONV2_MACoutF1_11  , In2_CONV2_MACoutF1_11  , In3_CONV2_MACoutF1_11  , In4_CONV2_MACoutF1_11  , Filter1BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F1_11 );


MUX5X1_13 F2_0 (In1_CONV2_MACoutF2_0  , In2_CONV2_MACoutF2_0  , In3_CONV2_MACoutF2_0  , In4_CONV2_MACoutF2_0  , Filter2BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F2_0 );
MUX5X1_13 F2_1 (In1_CONV2_MACoutF2_1  , In2_CONV2_MACoutF2_1  , In3_CONV2_MACoutF2_1  , In4_CONV2_MACoutF2_1  , Filter2BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F2_1 );
MUX5X1_13 F2_10 (In1_CONV2_MACoutF2_10  , In2_CONV2_MACoutF2_10  , In3_CONV2_MACoutF2_10  , In4_CONV2_MACoutF2_10  , Filter2BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F2_10 );
MUX5X1_13 F2_11 (In1_CONV2_MACoutF2_11  , In2_CONV2_MACoutF2_11  , In3_CONV2_MACoutF2_11  , In4_CONV2_MACoutF2_11  , Filter2BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F2_11 );


MUX5X1_13 F3_0 (In1_CONV2_MACoutF3_0  , In2_CONV2_MACoutF3_0  , In3_CONV2_MACoutF3_0  , In4_CONV2_MACoutF3_0  , Filter3BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F3_0 );
MUX5X1_13 F3_1 (In1_CONV2_MACoutF3_1  , In2_CONV2_MACoutF3_1  , In3_CONV2_MACoutF3_1  , In4_CONV2_MACoutF3_1  , Filter3BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F3_1 );
MUX5X1_13 F3_10 (In1_CONV2_MACoutF3_10  , In2_CONV2_MACoutF3_10  , In3_CONV2_MACoutF3_10  , In4_CONV2_MACoutF3_10  , Filter3BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F3_10 );
MUX5X1_13 F3_11 (In1_CONV2_MACoutF3_11  , In2_CONV2_MACoutF3_11  , In3_CONV2_MACoutF3_11  , In4_CONV2_MACoutF3_11  , Filter3BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F3_11 );


MUX5X1_13 F4_0 (In1_CONV2_MACoutF4_0  , In2_CONV2_MACoutF4_0  , In3_CONV2_MACoutF4_0  , In4_CONV2_MACoutF4_0  , Filter4BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F4_0 );
MUX5X1_13 F4_1 (In1_CONV2_MACoutF4_1  , In2_CONV2_MACoutF4_1  , In3_CONV2_MACoutF4_1  , In4_CONV2_MACoutF4_1  , Filter4BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F4_1 );
MUX5X1_13 F4_10 (In1_CONV2_MACoutF4_10  , In2_CONV2_MACoutF4_10  , In3_CONV2_MACoutF4_10  , In4_CONV2_MACoutF4_10  , Filter4BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F4_10 );
MUX5X1_13 F4_11 (In1_CONV2_MACoutF4_11  , In2_CONV2_MACoutF4_11  , In3_CONV2_MACoutF4_11  , In4_CONV2_MACoutF4_11  , Filter4BIASOUT, count_3bits, CONV2_Final_CONV2_MUXout_F4_11 );



wire[65:0] AdderF1Out0,AdderF1Out1,AdderF1Out10,AdderF1Out11;
wire[65:0] AdderF2Out0,AdderF2Out1,AdderF2Out10,AdderF2Out11;
wire[65:0] AdderF3Out0,AdderF3Out1,AdderF3Out10,AdderF3Out11;
wire[65:0] AdderF4Out0,AdderF4Out1,AdderF4Out10,AdderF4Out11;	



assign CONV2_MAC_start_Stage2 = (CONV2_counter >156)?1'b1 :1'b0; //(count_3bits >=2'b01) ?1'b1 :1'b0; //CONV2_MAC_end; 12*13 //156
assign  CONV2_MAC_end_Stage2=  (count_3bits >=63) ?1'b1 :1'b0; //5*13 65 64


AdderAcc_5 Adder_F1_0  (CONV2_Final_CONV2_MUXout_F1_0 , clk, AdderF1Out0  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F1_1  (CONV2_Final_CONV2_MUXout_F1_1 , clk, AdderF1Out1  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F1_10  (CONV2_Final_CONV2_MUXout_F1_10 , clk, AdderF1Out10  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F1_11  (CONV2_Final_CONV2_MUXout_F1_11 , clk, AdderF1Out11  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);

AdderAcc_5 Adder_F2_0  (CONV2_Final_CONV2_MUXout_F2_0 , clk, AdderF2Out0  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F2_1  (CONV2_Final_CONV2_MUXout_F2_1 , clk, AdderF2Out1  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F2_10  (CONV2_Final_CONV2_MUXout_F2_10 , clk, AdderF2Out10  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F2_11  (CONV2_Final_CONV2_MUXout_F2_11 , clk, AdderF2Out11  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);

AdderAcc_5 Adder_F3_0  (CONV2_Final_CONV2_MUXout_F3_0 , clk, AdderF3Out0  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F3_1  (CONV2_Final_CONV2_MUXout_F3_1 , clk, AdderF3Out1  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F3_10  (CONV2_Final_CONV2_MUXout_F3_10 , clk, AdderF3Out10  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F3_11  (CONV2_Final_CONV2_MUXout_F3_11 , clk, AdderF3Out11  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);

AdderAcc_5 Adder_F4_0  (CONV2_Final_CONV2_MUXout_F4_0 , clk, AdderF4Out0  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F4_1  (CONV2_Final_CONV2_MUXout_F4_1 , clk, AdderF4Out1  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F4_10  (CONV2_Final_CONV2_MUXout_F4_10 , clk, AdderF4Out10  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);
AdderAcc_5 Adder_F4_11  (CONV2_Final_CONV2_MUXout_F4_11 , clk, AdderF4Out11  , CONV2_MAC_start_Stage2, CONV2_MAC_end_Stage2, RST65);


wire[65:0] CONV2_RELU_F1out0,CONV2_RELU_F1out1,CONV2_RELU_F1out10,CONV2_RELU_F1out11;
wire[65:0] CONV2_RELU_F2out0,CONV2_RELU_F2out1,CONV2_RELU_F2out10,CONV2_RELU_F2out11;
wire[65:0] CONV2_RELU_F3out0,CONV2_RELU_F3out1,CONV2_RELU_F3out10,CONV2_RELU_F3out11;
wire[65:0] CONV2_RELU_F4out0,CONV2_RELU_F4out1,CONV2_RELU_F4out10,CONV2_RELU_F4out11;


RELU Conv2RELU_F1_0 (AdderF1Out0  , clk , CONV2_RELU_F1out0 );
RELU Conv2RELU_F1_1 (AdderF1Out1  , clk , CONV2_RELU_F1out1 );
RELU Conv2RELU_F1_10 (AdderF1Out10  , clk , CONV2_RELU_F1out10 );
RELU Conv2RELU_F1_11 (AdderF1Out11  , clk , CONV2_RELU_F1out11 );

RELU Conv2RELU_F2_0 (AdderF2Out0  , clk , CONV2_RELU_F2out0 );
RELU Conv2RELU_F2_1 (AdderF2Out1  , clk , CONV2_RELU_F2out1 );
RELU Conv2RELU_F2_10 (AdderF2Out10  , clk , CONV2_RELU_F2out10 );
RELU Conv2RELU_F2_11 (AdderF2Out11  , clk , CONV2_RELU_F2out11 );

RELU Conv2RELU_F3_0 (AdderF3Out0  , clk , CONV2_RELU_F3out0 );
RELU Conv2RELU_F3_1 (AdderF3Out1  , clk , CONV2_RELU_F3out1 );
RELU Conv2RELU_F3_10 (AdderF3Out10  , clk , CONV2_RELU_F3out10 );
RELU Conv2RELU_F3_11 (AdderF3Out11  , clk , CONV2_RELU_F3out11 );

RELU Conv2RELU_F4_0 (AdderF4Out0  , clk , CONV2_RELU_F4out0 );
RELU Conv2RELU_F4_1 (AdderF4Out1  , clk , CONV2_RELU_F4out1 );
RELU Conv2RELU_F4_10 (AdderF4Out10  , clk , CONV2_RELU_F4out10 );
RELU Conv2RELU_F4_11 (AdderF4Out11  , clk , CONV2_RELU_F4out11 );



assign LayerStartStage2 = (CONV2_counter >154)?1'b1 :1'b0; //156 jjjj

reg Stage2_xwrite_1 , Stage2_xwrite_2, Stage2_xwrite_3, Stage2_xwrite_4, Stage2_xwrite_5;
reg Stage2_xwrite_6 , Stage2_xwrite_7, Stage2_xwrite_8, Stage2_xwrite_9, Stage2_xwrite_10;
reg  Stage2_xwrite_11, Stage2_xwrite_12, Stage2_xwrite_13, Stage2_xwrite_14, Stage2_xwrite_15;
reg Stage2_xwrite_16 , Stage2_xwrite_17, Stage2_xwrite_18, Stage2_xwrite_19, Stage2_xwrite_20;
reg Stage2_xwrite_21 , Stage2_xwrite_22 , Stage2_xwrite_23, Stage2_xwrite_24, Stage2_xwrite_25;



always @ (posedge clk)
begin

if (bigaddress ==  0) begin resetTheCounter <= 1;

Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;

end

else if (bigaddress ==   221) begin resetTheCounter <= 1; //
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   223) begin resetTheCounter <= 0; //
Stage2_xwrite_1 <= 1; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end

else if (bigaddress ==   443) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   444) begin resetTheCounter <= 0; //444
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 1; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end

else if (bigaddress ==   665) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end
else if (bigaddress ==   666) begin resetTheCounter <= 0; //666
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 1; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end

else if (bigaddress ==   887) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   888) begin resetTheCounter <= 0;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 1; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   1109 ) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   1110 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 1;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   1331) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   1332 ) begin resetTheCounter <= 0; //
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 1; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   1553) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   1554 ) begin resetTheCounter <= 0; //
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 1; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   1775) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   1776 ) begin resetTheCounter <= 0; //
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 1; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   1997) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   1998 ) begin resetTheCounter <= 0; //
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 1; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end

else if (bigaddress ==   2219) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   2220 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 1;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   2441) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   2442 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 1; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   2663) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   2664 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 1; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   2885) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   2886 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 1; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   3107) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   3108 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 1; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   3329) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   3330 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 1;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   3551 ) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   3552  ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 1; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   3773) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   3774 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 1; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   3995) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   3996 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 1; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end



else if (bigaddress ==   4217 ) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   4218  ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 1; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0; 
end


else if (bigaddress ==   4439) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==  4440  ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 1;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end

else if (bigaddress ==   4661) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   4662 ) begin resetTheCounter <= 0; //
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 1; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end

else if (bigaddress ==   4883 ) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   4884  ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 1; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   5105) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   5106 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 1; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   5327) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   5328 ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 1; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   5549 ) begin resetTheCounter <= 1;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end


else if (bigaddress ==   5550  ) begin resetTheCounter <= 0;//
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 1;
end


else begin resetTheCounter <= 0;
Stage2_xwrite_1 <= 0; Stage2_xwrite_2 <= 0; Stage2_xwrite_3 <= 0; Stage2_xwrite_4 <= 0; Stage2_xwrite_5 <= 0;
Stage2_xwrite_6 <= 0; Stage2_xwrite_7<= 0; Stage2_xwrite_8 <= 0; Stage2_xwrite_9 <= 0; Stage2_xwrite_10 <= 0;
Stage2_xwrite_11 <= 0; Stage2_xwrite_12 <= 0; Stage2_xwrite_13 <= 0; Stage2_xwrite_14 <= 0; Stage2_xwrite_15 <= 0;
Stage2_xwrite_16 <= 0; Stage2_xwrite_17 <= 0; Stage2_xwrite_18 <= 0; Stage2_xwrite_19 <= 0; Stage2_xwrite_20 <= 0;
Stage2_xwrite_21 <= 0; Stage2_xwrite_22 <= 0; Stage2_xwrite_23 <= 0; Stage2_xwrite_24 <= 0; Stage2_xwrite_25 <= 0;
end
end



OneRegisterOut RAMFilter1Combined0  (clk, Stage2_xwrite_1, CONV2_RELU_F1out0 , LastRamOutF1_0 );
OneRegisterOut RAMFilter1Combined1  (clk, Stage2_xwrite_1, CONV2_RELU_F1out1 , LastRamOutF1_1 );
OneRegisterOut RAMFilter1Combined2  (clk, Stage2_xwrite_2, CONV2_RELU_F1out0 , LastRamOutF1_2 );
OneRegisterOut RAMFilter1Combined3  (clk, Stage2_xwrite_2, CONV2_RELU_F1out1 , LastRamOutF1_3 );
OneRegisterOut RAMFilter1Combined4  (clk, Stage2_xwrite_3, CONV2_RELU_F1out0 , LastRamOutF1_4 );
OneRegisterOut RAMFilter1Combined5  (clk, Stage2_xwrite_3, CONV2_RELU_F1out1 , LastRamOutF1_5 );
OneRegisterOut RAMFilter1Combined6  (clk, Stage2_xwrite_4, CONV2_RELU_F1out0 , LastRamOutF1_6 );
OneRegisterOut RAMFilter1Combined7  (clk, Stage2_xwrite_4, CONV2_RELU_F1out1 , LastRamOutF1_7 );
OneRegisterOut RAMFilter1Combined8  (clk, Stage2_xwrite_5, CONV2_RELU_F1out0 , LastRamOutF1_8 );
OneRegisterOut RAMFilter1Combined9  (clk, Stage2_xwrite_5, CONV2_RELU_F1out1 , LastRamOutF1_9 );


OneRegisterOut RAMFilter1Combined10  (clk, Stage2_xwrite_1, CONV2_RELU_F1out10 , LastRamOutF1_10 );
OneRegisterOut RAMFilter1Combined11  (clk, Stage2_xwrite_1, CONV2_RELU_F1out11 , LastRamOutF1_11 );
OneRegisterOut RAMFilter1Combined12  (clk, Stage2_xwrite_2, CONV2_RELU_F1out10 , LastRamOutF1_12 );
OneRegisterOut RAMFilter1Combined13  (clk, Stage2_xwrite_2, CONV2_RELU_F1out11 , LastRamOutF1_13 );
OneRegisterOut RAMFilter1Combined14  (clk, Stage2_xwrite_3, CONV2_RELU_F1out10 , LastRamOutF1_14 );
OneRegisterOut RAMFilter1Combined15  (clk, Stage2_xwrite_3, CONV2_RELU_F1out11 , LastRamOutF1_15 );
OneRegisterOut RAMFilter1Combined16  (clk, Stage2_xwrite_4, CONV2_RELU_F1out10 , LastRamOutF1_16 );
OneRegisterOut RAMFilter1Combined17  (clk, Stage2_xwrite_4, CONV2_RELU_F1out11 , LastRamOutF1_17 );
OneRegisterOut RAMFilter1Combined18  (clk, Stage2_xwrite_5, CONV2_RELU_F1out10 , LastRamOutF1_18 );
OneRegisterOut RAMFilter1Combined19  (clk, Stage2_xwrite_5, CONV2_RELU_F1out11 , LastRamOutF1_19 );



OneRegisterOut RAMFilter1Combined20  (clk, Stage2_xwrite_6, CONV2_RELU_F1out0 , LastRamOutF1_20 );
OneRegisterOut RAMFilter1Combined21  (clk, Stage2_xwrite_6, CONV2_RELU_F1out1 , LastRamOutF1_21 );
OneRegisterOut RAMFilter1Combined22  (clk, Stage2_xwrite_7, CONV2_RELU_F1out0 , LastRamOutF1_22 );
OneRegisterOut RAMFilter1Combined23  (clk, Stage2_xwrite_7, CONV2_RELU_F1out1 , LastRamOutF1_23 );
OneRegisterOut RAMFilter1Combined24  (clk, Stage2_xwrite_8, CONV2_RELU_F1out0 , LastRamOutF1_24 );
OneRegisterOut RAMFilter1Combined25  (clk, Stage2_xwrite_8, CONV2_RELU_F1out1 , LastRamOutF1_25 );
OneRegisterOut RAMFilter1Combined26  (clk, Stage2_xwrite_9, CONV2_RELU_F1out0 , LastRamOutF1_26 );
OneRegisterOut RAMFilter1Combined27  (clk, Stage2_xwrite_9, CONV2_RELU_F1out1 , LastRamOutF1_27 );
OneRegisterOut RAMFilter1Combined28  (clk, Stage2_xwrite_10, CONV2_RELU_F1out0 , LastRamOutF1_28 );
OneRegisterOut RAMFilter1Combined29  (clk, Stage2_xwrite_10, CONV2_RELU_F1out1 , LastRamOutF1_29 );


OneRegisterOut RAMFilter1Combined30  (clk, Stage2_xwrite_6, CONV2_RELU_F1out10 , LastRamOutF1_30 );
OneRegisterOut RAMFilter1Combined31  (clk, Stage2_xwrite_6, CONV2_RELU_F1out11 , LastRamOutF1_31 );
OneRegisterOut RAMFilter1Combined32  (clk, Stage2_xwrite_7, CONV2_RELU_F1out10 , LastRamOutF1_32 );
OneRegisterOut RAMFilter1Combined33  (clk, Stage2_xwrite_7, CONV2_RELU_F1out11 , LastRamOutF1_33 );
OneRegisterOut RAMFilter1Combined34  (clk, Stage2_xwrite_8, CONV2_RELU_F1out10 , LastRamOutF1_34 );
OneRegisterOut RAMFilter1Combined35  (clk, Stage2_xwrite_8, CONV2_RELU_F1out11 , LastRamOutF1_35 );
OneRegisterOut RAMFilter1Combined36  (clk, Stage2_xwrite_9, CONV2_RELU_F1out10 , LastRamOutF1_36 );
OneRegisterOut RAMFilter1Combined37  (clk, Stage2_xwrite_9, CONV2_RELU_F1out11 , LastRamOutF1_37 );
OneRegisterOut RAMFilter1Combined38  (clk, Stage2_xwrite_10, CONV2_RELU_F1out10 , LastRamOutF1_38 );
OneRegisterOut RAMFilter1Combined39  (clk, Stage2_xwrite_10, CONV2_RELU_F1out11 , LastRamOutF1_39 );



OneRegisterOut RAMFilter1Combined40  (clk, Stage2_xwrite_11, CONV2_RELU_F1out0 , LastRamOutF1_40 );
OneRegisterOut RAMFilter1Combined41  (clk, Stage2_xwrite_11, CONV2_RELU_F1out1 , LastRamOutF1_41 );
OneRegisterOut RAMFilter1Combined42  (clk, Stage2_xwrite_12, CONV2_RELU_F1out0 , LastRamOutF1_42 );
OneRegisterOut RAMFilter1Combined43  (clk, Stage2_xwrite_12, CONV2_RELU_F1out1 , LastRamOutF1_43 );
OneRegisterOut RAMFilter1Combined44  (clk, Stage2_xwrite_13, CONV2_RELU_F1out0 , LastRamOutF1_44 );
OneRegisterOut RAMFilter1Combined45  (clk, Stage2_xwrite_13, CONV2_RELU_F1out1 , LastRamOutF1_45 );
OneRegisterOut RAMFilter1Combined46  (clk, Stage2_xwrite_14, CONV2_RELU_F1out0 , LastRamOutF1_46 );
OneRegisterOut RAMFilter1Combined47  (clk, Stage2_xwrite_14, CONV2_RELU_F1out1 , LastRamOutF1_47 );
OneRegisterOut RAMFilter1Combined48  (clk, Stage2_xwrite_15, CONV2_RELU_F1out0 , LastRamOutF1_48 );
OneRegisterOut RAMFilter1Combined49  (clk, Stage2_xwrite_15, CONV2_RELU_F1out1 , LastRamOutF1_49 );


OneRegisterOut RAMFilter1Combined50  (clk, Stage2_xwrite_11, CONV2_RELU_F1out10 , LastRamOutF1_50 );
OneRegisterOut RAMFilter1Combined51  (clk, Stage2_xwrite_11, CONV2_RELU_F1out11 , LastRamOutF1_51 );
OneRegisterOut RAMFilter1Combined52  (clk, Stage2_xwrite_12, CONV2_RELU_F1out10 , LastRamOutF1_52 );
OneRegisterOut RAMFilter1Combined53  (clk, Stage2_xwrite_12, CONV2_RELU_F1out11 , LastRamOutF1_53 );
OneRegisterOut RAMFilter1Combined54  (clk, Stage2_xwrite_13, CONV2_RELU_F1out10 , LastRamOutF1_54 );
OneRegisterOut RAMFilter1Combined55  (clk, Stage2_xwrite_13, CONV2_RELU_F1out11 , LastRamOutF1_55 );
OneRegisterOut RAMFilter1Combined56  (clk, Stage2_xwrite_14, CONV2_RELU_F1out10 , LastRamOutF1_56 );
OneRegisterOut RAMFilter1Combined57  (clk, Stage2_xwrite_14, CONV2_RELU_F1out11 , LastRamOutF1_57 );
OneRegisterOut RAMFilter1Combined58  (clk, Stage2_xwrite_15, CONV2_RELU_F1out10 , LastRamOutF1_58 );
OneRegisterOut RAMFilter1Combined59  (clk, Stage2_xwrite_15, CONV2_RELU_F1out11 , LastRamOutF1_59 );




OneRegisterOut RAMFilter1Combined60  (clk, Stage2_xwrite_16, CONV2_RELU_F1out0 , LastRamOutF1_60 );
OneRegisterOut RAMFilter1Combined61  (clk, Stage2_xwrite_16, CONV2_RELU_F1out1 , LastRamOutF1_61 );
OneRegisterOut RAMFilter1Combined62  (clk, Stage2_xwrite_17, CONV2_RELU_F1out0 , LastRamOutF1_62 );
OneRegisterOut RAMFilter1Combined63  (clk, Stage2_xwrite_17, CONV2_RELU_F1out1 , LastRamOutF1_63 );
OneRegisterOut RAMFilter1Combined64  (clk, Stage2_xwrite_18, CONV2_RELU_F1out0 , LastRamOutF1_64 );
OneRegisterOut RAMFilter1Combined65  (clk, Stage2_xwrite_18, CONV2_RELU_F1out1 , LastRamOutF1_65 );
OneRegisterOut RAMFilter1Combined66  (clk, Stage2_xwrite_19, CONV2_RELU_F1out0 , LastRamOutF1_66 );
OneRegisterOut RAMFilter1Combined67  (clk, Stage2_xwrite_19, CONV2_RELU_F1out1 , LastRamOutF1_67 );
OneRegisterOut RAMFilter1Combined68  (clk, Stage2_xwrite_20, CONV2_RELU_F1out0 , LastRamOutF1_68 );
OneRegisterOut RAMFilter1Combined69  (clk, Stage2_xwrite_20, CONV2_RELU_F1out1 , LastRamOutF1_69 );


OneRegisterOut RAMFilter1Combined70  (clk, Stage2_xwrite_16, CONV2_RELU_F1out10 , LastRamOutF1_70 );
OneRegisterOut RAMFilter1Combined71  (clk, Stage2_xwrite_16, CONV2_RELU_F1out11 , LastRamOutF1_71 );
OneRegisterOut RAMFilter1Combined72  (clk, Stage2_xwrite_17, CONV2_RELU_F1out10 , LastRamOutF1_72 );
OneRegisterOut RAMFilter1Combined73  (clk, Stage2_xwrite_17, CONV2_RELU_F1out11 , LastRamOutF1_73 );
OneRegisterOut RAMFilter1Combined74  (clk, Stage2_xwrite_18, CONV2_RELU_F1out10 , LastRamOutF1_74 );
OneRegisterOut RAMFilter1Combined75  (clk, Stage2_xwrite_18, CONV2_RELU_F1out11 , LastRamOutF1_75 );
OneRegisterOut RAMFilter1Combined76  (clk, Stage2_xwrite_19, CONV2_RELU_F1out10 , LastRamOutF1_76 );
OneRegisterOut RAMFilter1Combined77  (clk, Stage2_xwrite_19, CONV2_RELU_F1out11 , LastRamOutF1_77 );
OneRegisterOut RAMFilter1Combined78  (clk, Stage2_xwrite_20, CONV2_RELU_F1out10 , LastRamOutF1_78 );
OneRegisterOut RAMFilter1Combined79  (clk, Stage2_xwrite_20, CONV2_RELU_F1out11 , LastRamOutF1_79 );



OneRegisterOut RAMFilter1Combined80  (clk, Stage2_xwrite_21, CONV2_RELU_F1out0 , LastRamOutF1_80 );
OneRegisterOut RAMFilter1Combined81  (clk, Stage2_xwrite_21, CONV2_RELU_F1out1 , LastRamOutF1_81 );
OneRegisterOut RAMFilter1Combined82  (clk, Stage2_xwrite_22, CONV2_RELU_F1out0 , LastRamOutF1_82 );
OneRegisterOut RAMFilter1Combined83  (clk, Stage2_xwrite_22, CONV2_RELU_F1out1 , LastRamOutF1_83 );
OneRegisterOut RAMFilter1Combined84  (clk, Stage2_xwrite_23, CONV2_RELU_F1out0 , LastRamOutF1_84 );
OneRegisterOut RAMFilter1Combined85  (clk, Stage2_xwrite_23, CONV2_RELU_F1out1 , LastRamOutF1_85 );
OneRegisterOut RAMFilter1Combined86  (clk, Stage2_xwrite_24, CONV2_RELU_F1out0 , LastRamOutF1_86 );
OneRegisterOut RAMFilter1Combined87  (clk, Stage2_xwrite_24, CONV2_RELU_F1out1 , LastRamOutF1_87 );
OneRegisterOut RAMFilter1Combined88  (clk, Stage2_xwrite_25, CONV2_RELU_F1out0 , LastRamOutF1_88 );
OneRegisterOut RAMFilter1Combined89  (clk, Stage2_xwrite_25, CONV2_RELU_F1out1 , LastRamOutF1_89 );


OneRegisterOut RAMFilter1Combined90  (clk, Stage2_xwrite_21, CONV2_RELU_F1out10 , LastRamOutF1_90 );
OneRegisterOut RAMFilter1Combined91  (clk, Stage2_xwrite_21, CONV2_RELU_F1out11 , LastRamOutF1_91 );
OneRegisterOut RAMFilter1Combined92  (clk, Stage2_xwrite_22, CONV2_RELU_F1out10 , LastRamOutF1_92 );
OneRegisterOut RAMFilter1Combined93  (clk, Stage2_xwrite_22, CONV2_RELU_F1out11 , LastRamOutF1_93 );
OneRegisterOut RAMFilter1Combined94  (clk, Stage2_xwrite_23, CONV2_RELU_F1out10 , LastRamOutF1_94 );
OneRegisterOut RAMFilter1Combined95  (clk, Stage2_xwrite_23, CONV2_RELU_F1out11 , LastRamOutF1_95 );
OneRegisterOut RAMFilter1Combined96  (clk, Stage2_xwrite_24, CONV2_RELU_F1out10 , LastRamOutF1_96 );
OneRegisterOut RAMFilter1Combined97  (clk, Stage2_xwrite_24, CONV2_RELU_F1out11 , LastRamOutF1_97 );
OneRegisterOut RAMFilter1Combined98  (clk, Stage2_xwrite_25, CONV2_RELU_F1out10 , LastRamOutF1_98 );
OneRegisterOut RAMFilter1Combined99  (clk, Stage2_xwrite_25, CONV2_RELU_F1out11 , LastRamOutF1_99 );


///



OneRegisterOut RAMFilter2Combined0  (clk, Stage2_xwrite_1, CONV2_RELU_F2out0 , LastRamOutF2_0 );
OneRegisterOut RAMFilter2Combined1  (clk, Stage2_xwrite_1, CONV2_RELU_F2out1 , LastRamOutF2_1 );
OneRegisterOut RAMFilter2Combined2  (clk, Stage2_xwrite_2, CONV2_RELU_F2out0 , LastRamOutF2_2 );
OneRegisterOut RAMFilter2Combined3  (clk, Stage2_xwrite_2, CONV2_RELU_F2out1 , LastRamOutF2_3 );
OneRegisterOut RAMFilter2Combined4  (clk, Stage2_xwrite_3, CONV2_RELU_F2out0 , LastRamOutF2_4 );
OneRegisterOut RAMFilter2Combined5  (clk, Stage2_xwrite_3, CONV2_RELU_F2out1 , LastRamOutF2_5 );
OneRegisterOut RAMFilter2Combined6  (clk, Stage2_xwrite_4, CONV2_RELU_F2out0 , LastRamOutF2_6 );
OneRegisterOut RAMFilter2Combined7  (clk, Stage2_xwrite_4, CONV2_RELU_F2out1 , LastRamOutF2_7 );
OneRegisterOut RAMFilter2Combined8  (clk, Stage2_xwrite_5, CONV2_RELU_F2out0 , LastRamOutF2_8 );
OneRegisterOut RAMFilter2Combined9  (clk, Stage2_xwrite_5, CONV2_RELU_F2out1 , LastRamOutF2_9 );

OneRegisterOut RAMFilter2Combined10  (clk, Stage2_xwrite_1, CONV2_RELU_F2out10 , LastRamOutF2_10 );
OneRegisterOut RAMFilter2Combined11  (clk, Stage2_xwrite_1, CONV2_RELU_F2out11 , LastRamOutF2_11 );
OneRegisterOut RAMFilter2Combined12  (clk, Stage2_xwrite_2, CONV2_RELU_F2out10 , LastRamOutF2_12 );
OneRegisterOut RAMFilter2Combined13  (clk, Stage2_xwrite_2, CONV2_RELU_F2out11 , LastRamOutF2_13 );
OneRegisterOut RAMFilter2Combined14  (clk, Stage2_xwrite_3, CONV2_RELU_F2out10 , LastRamOutF2_14 );
OneRegisterOut RAMFilter2Combined15  (clk, Stage2_xwrite_3, CONV2_RELU_F2out11 , LastRamOutF2_15 );
OneRegisterOut RAMFilter2Combined16  (clk, Stage2_xwrite_4, CONV2_RELU_F2out10 , LastRamOutF2_16 );
OneRegisterOut RAMFilter2Combined17  (clk, Stage2_xwrite_4, CONV2_RELU_F2out11 , LastRamOutF2_17 );
OneRegisterOut RAMFilter2Combined18  (clk, Stage2_xwrite_5, CONV2_RELU_F2out10 , LastRamOutF2_18 );
OneRegisterOut RAMFilter2Combined19  (clk, Stage2_xwrite_5, CONV2_RELU_F2out11 , LastRamOutF2_19 );

OneRegisterOut RAMFilter2Combined20  (clk, Stage2_xwrite_6, CONV2_RELU_F2out0 , LastRamOutF2_20 );
OneRegisterOut RAMFilter2Combined21  (clk, Stage2_xwrite_6, CONV2_RELU_F2out1 , LastRamOutF2_21 );
OneRegisterOut RAMFilter2Combined22  (clk, Stage2_xwrite_7, CONV2_RELU_F2out0 , LastRamOutF2_22 );
OneRegisterOut RAMFilter2Combined23  (clk, Stage2_xwrite_7, CONV2_RELU_F2out1 , LastRamOutF2_23 );
OneRegisterOut RAMFilter2Combined24  (clk, Stage2_xwrite_8, CONV2_RELU_F2out0 , LastRamOutF2_24 );
OneRegisterOut RAMFilter2Combined25  (clk, Stage2_xwrite_8, CONV2_RELU_F2out1 , LastRamOutF2_25 );
OneRegisterOut RAMFilter2Combined26  (clk, Stage2_xwrite_9, CONV2_RELU_F2out0 , LastRamOutF2_26 );
OneRegisterOut RAMFilter2Combined27  (clk, Stage2_xwrite_9, CONV2_RELU_F2out1 , LastRamOutF2_27 );
OneRegisterOut RAMFilter2Combined28  (clk, Stage2_xwrite_10, CONV2_RELU_F2out0 , LastRamOutF2_28 );
OneRegisterOut RAMFilter2Combined29  (clk, Stage2_xwrite_10, CONV2_RELU_F2out1 , LastRamOutF2_29 );

OneRegisterOut RAMFilter2Combined30  (clk, Stage2_xwrite_6, CONV2_RELU_F2out10 , LastRamOutF2_30 );
OneRegisterOut RAMFilter2Combined31  (clk, Stage2_xwrite_6, CONV2_RELU_F2out11 , LastRamOutF2_31 );
OneRegisterOut RAMFilter2Combined32  (clk, Stage2_xwrite_7, CONV2_RELU_F2out10 , LastRamOutF2_32 );
OneRegisterOut RAMFilter2Combined33  (clk, Stage2_xwrite_7, CONV2_RELU_F2out11 , LastRamOutF2_33 );
OneRegisterOut RAMFilter2Combined34  (clk, Stage2_xwrite_8, CONV2_RELU_F2out10 , LastRamOutF2_34 );
OneRegisterOut RAMFilter2Combined35  (clk, Stage2_xwrite_8, CONV2_RELU_F2out11 , LastRamOutF2_35 );
OneRegisterOut RAMFilter2Combined36  (clk, Stage2_xwrite_9, CONV2_RELU_F2out10 , LastRamOutF2_36 );
OneRegisterOut RAMFilter2Combined37  (clk, Stage2_xwrite_9, CONV2_RELU_F2out11 , LastRamOutF2_37 );
OneRegisterOut RAMFilter2Combined38  (clk, Stage2_xwrite_10, CONV2_RELU_F2out10 , LastRamOutF2_38 );
OneRegisterOut RAMFilter2Combined39  (clk, Stage2_xwrite_10, CONV2_RELU_F2out11 , LastRamOutF2_39 );

OneRegisterOut RAMFilter2Combined40  (clk, Stage2_xwrite_11, CONV2_RELU_F2out0 , LastRamOutF2_40 );
OneRegisterOut RAMFilter2Combined41  (clk, Stage2_xwrite_11, CONV2_RELU_F2out1 , LastRamOutF2_41 );
OneRegisterOut RAMFilter2Combined42  (clk, Stage2_xwrite_12, CONV2_RELU_F2out0 , LastRamOutF2_42 );
OneRegisterOut RAMFilter2Combined43  (clk, Stage2_xwrite_12, CONV2_RELU_F2out1 , LastRamOutF2_43 );
OneRegisterOut RAMFilter2Combined44  (clk, Stage2_xwrite_13, CONV2_RELU_F2out0 , LastRamOutF2_44 );
OneRegisterOut RAMFilter2Combined45  (clk, Stage2_xwrite_13, CONV2_RELU_F2out1 , LastRamOutF2_45 );
OneRegisterOut RAMFilter2Combined46  (clk, Stage2_xwrite_14, CONV2_RELU_F2out0 , LastRamOutF2_46 );
OneRegisterOut RAMFilter2Combined47  (clk, Stage2_xwrite_14, CONV2_RELU_F2out1 , LastRamOutF2_47 );
OneRegisterOut RAMFilter2Combined48  (clk, Stage2_xwrite_15, CONV2_RELU_F2out0 , LastRamOutF2_48 );
OneRegisterOut RAMFilter2Combined49  (clk, Stage2_xwrite_15, CONV2_RELU_F2out1 , LastRamOutF2_49 );

OneRegisterOut RAMFilter2Combined50  (clk, Stage2_xwrite_11, CONV2_RELU_F2out10 , LastRamOutF2_50 );
OneRegisterOut RAMFilter2Combined51  (clk, Stage2_xwrite_11, CONV2_RELU_F2out11 , LastRamOutF2_51 );
OneRegisterOut RAMFilter2Combined52  (clk, Stage2_xwrite_12, CONV2_RELU_F2out10 , LastRamOutF2_52 );
OneRegisterOut RAMFilter2Combined53  (clk, Stage2_xwrite_12, CONV2_RELU_F2out11 , LastRamOutF2_53 );
OneRegisterOut RAMFilter2Combined54  (clk, Stage2_xwrite_13, CONV2_RELU_F2out10 , LastRamOutF2_54 );
OneRegisterOut RAMFilter2Combined55  (clk, Stage2_xwrite_13, CONV2_RELU_F2out11 , LastRamOutF2_55 );
OneRegisterOut RAMFilter2Combined56  (clk, Stage2_xwrite_14, CONV2_RELU_F2out10 , LastRamOutF2_56 );
OneRegisterOut RAMFilter2Combined57  (clk, Stage2_xwrite_14, CONV2_RELU_F2out11 , LastRamOutF2_57 );
OneRegisterOut RAMFilter2Combined58  (clk, Stage2_xwrite_15, CONV2_RELU_F2out10 , LastRamOutF2_58 );
OneRegisterOut RAMFilter2Combined59  (clk, Stage2_xwrite_15, CONV2_RELU_F2out11 , LastRamOutF2_59 );

OneRegisterOut RAMFilter2Combined60  (clk, Stage2_xwrite_16, CONV2_RELU_F2out0 , LastRamOutF2_60 );
OneRegisterOut RAMFilter2Combined61  (clk, Stage2_xwrite_16, CONV2_RELU_F2out1 , LastRamOutF2_61 );
OneRegisterOut RAMFilter2Combined62  (clk, Stage2_xwrite_17, CONV2_RELU_F2out0 , LastRamOutF2_62 );
OneRegisterOut RAMFilter2Combined63  (clk, Stage2_xwrite_17, CONV2_RELU_F2out1 , LastRamOutF2_63 );
OneRegisterOut RAMFilter2Combined64  (clk, Stage2_xwrite_18, CONV2_RELU_F2out0 , LastRamOutF2_64 );
OneRegisterOut RAMFilter2Combined65  (clk, Stage2_xwrite_18, CONV2_RELU_F2out1 , LastRamOutF2_65 );
OneRegisterOut RAMFilter2Combined66  (clk, Stage2_xwrite_19, CONV2_RELU_F2out0 , LastRamOutF2_66 );
OneRegisterOut RAMFilter2Combined67  (clk, Stage2_xwrite_19, CONV2_RELU_F2out1 , LastRamOutF2_67 );
OneRegisterOut RAMFilter2Combined68  (clk, Stage2_xwrite_20, CONV2_RELU_F2out0 , LastRamOutF2_68 );
OneRegisterOut RAMFilter2Combined69  (clk, Stage2_xwrite_20, CONV2_RELU_F2out1 , LastRamOutF2_69 );

OneRegisterOut RAMFilter2Combined70  (clk, Stage2_xwrite_16, CONV2_RELU_F2out10 , LastRamOutF2_70 );
OneRegisterOut RAMFilter2Combined71  (clk, Stage2_xwrite_16, CONV2_RELU_F2out11 , LastRamOutF2_71 );
OneRegisterOut RAMFilter2Combined72  (clk, Stage2_xwrite_17, CONV2_RELU_F2out10 , LastRamOutF2_72 );
OneRegisterOut RAMFilter2Combined73  (clk, Stage2_xwrite_17, CONV2_RELU_F2out11 , LastRamOutF2_73 );
OneRegisterOut RAMFilter2Combined74  (clk, Stage2_xwrite_18, CONV2_RELU_F2out10 , LastRamOutF2_74 );
OneRegisterOut RAMFilter2Combined75  (clk, Stage2_xwrite_18, CONV2_RELU_F2out11 , LastRamOutF2_75 );
OneRegisterOut RAMFilter2Combined76  (clk, Stage2_xwrite_19, CONV2_RELU_F2out10 , LastRamOutF2_76 );
OneRegisterOut RAMFilter2Combined77  (clk, Stage2_xwrite_19, CONV2_RELU_F2out11 , LastRamOutF2_77 );
OneRegisterOut RAMFilter2Combined78  (clk, Stage2_xwrite_20, CONV2_RELU_F2out10 , LastRamOutF2_78 );
OneRegisterOut RAMFilter2Combined79  (clk, Stage2_xwrite_20, CONV2_RELU_F2out11 , LastRamOutF2_79 );

OneRegisterOut RAMFilter2Combined80  (clk, Stage2_xwrite_21, CONV2_RELU_F2out0 , LastRamOutF2_80 );
OneRegisterOut RAMFilter2Combined81  (clk, Stage2_xwrite_21, CONV2_RELU_F2out1 , LastRamOutF2_81 );
OneRegisterOut RAMFilter2Combined82  (clk, Stage2_xwrite_22, CONV2_RELU_F2out0 , LastRamOutF2_82 );
OneRegisterOut RAMFilter2Combined83  (clk, Stage2_xwrite_22, CONV2_RELU_F2out1 , LastRamOutF2_83 );
OneRegisterOut RAMFilter2Combined84  (clk, Stage2_xwrite_23, CONV2_RELU_F2out0 , LastRamOutF2_84 );
OneRegisterOut RAMFilter2Combined85  (clk, Stage2_xwrite_23, CONV2_RELU_F2out1 , LastRamOutF2_85 );
OneRegisterOut RAMFilter2Combined86  (clk, Stage2_xwrite_24, CONV2_RELU_F2out0 , LastRamOutF2_86 );
OneRegisterOut RAMFilter2Combined87  (clk, Stage2_xwrite_24, CONV2_RELU_F2out1 , LastRamOutF2_87 );
OneRegisterOut RAMFilter2Combined88  (clk, Stage2_xwrite_25, CONV2_RELU_F2out0 , LastRamOutF2_88 );
OneRegisterOut RAMFilter2Combined89  (clk, Stage2_xwrite_25, CONV2_RELU_F2out1 , LastRamOutF2_89 );

OneRegisterOut RAMFilter2Combined90  (clk, Stage2_xwrite_21, CONV2_RELU_F2out10 , LastRamOutF2_90 );
OneRegisterOut RAMFilter2Combined91  (clk, Stage2_xwrite_21, CONV2_RELU_F2out11 , LastRamOutF2_91 );
OneRegisterOut RAMFilter2Combined92  (clk, Stage2_xwrite_22, CONV2_RELU_F2out10 , LastRamOutF2_92 );
OneRegisterOut RAMFilter2Combined93  (clk, Stage2_xwrite_22, CONV2_RELU_F2out11 , LastRamOutF2_93 );
OneRegisterOut RAMFilter2Combined94  (clk, Stage2_xwrite_23, CONV2_RELU_F2out10 , LastRamOutF2_94 );
OneRegisterOut RAMFilter2Combined95  (clk, Stage2_xwrite_23, CONV2_RELU_F2out11 , LastRamOutF2_95 );
OneRegisterOut RAMFilter2Combined96  (clk, Stage2_xwrite_24, CONV2_RELU_F2out10 , LastRamOutF2_96 );
OneRegisterOut RAMFilter2Combined97  (clk, Stage2_xwrite_24, CONV2_RELU_F2out11 , LastRamOutF2_97 );
OneRegisterOut RAMFilter2Combined98  (clk, Stage2_xwrite_25, CONV2_RELU_F2out10 , LastRamOutF2_98 );
OneRegisterOut RAMFilter2Combined99  (clk, Stage2_xwrite_25, CONV2_RELU_F2out11 , LastRamOutF2_99 );

///



OneRegisterOut RAMFilter3Combined0  (clk, Stage2_xwrite_1, CONV2_RELU_F3out0 , LastRamOutF3_0 );
OneRegisterOut RAMFilter3Combined1  (clk, Stage2_xwrite_1, CONV2_RELU_F3out1 , LastRamOutF3_1 );
OneRegisterOut RAMFilter3Combined2  (clk, Stage2_xwrite_2, CONV2_RELU_F3out0 , LastRamOutF3_2 );
OneRegisterOut RAMFilter3Combined3  (clk, Stage2_xwrite_2, CONV2_RELU_F3out1 , LastRamOutF3_3 );
OneRegisterOut RAMFilter3Combined4  (clk, Stage2_xwrite_3, CONV2_RELU_F3out0 , LastRamOutF3_4 );
OneRegisterOut RAMFilter3Combined5  (clk, Stage2_xwrite_3, CONV2_RELU_F3out1 , LastRamOutF3_5 );
OneRegisterOut RAMFilter3Combined6  (clk, Stage2_xwrite_4, CONV2_RELU_F3out0 , LastRamOutF3_6 );
OneRegisterOut RAMFilter3Combined7  (clk, Stage2_xwrite_4, CONV2_RELU_F3out1 , LastRamOutF3_7 );
OneRegisterOut RAMFilter3Combined8  (clk, Stage2_xwrite_5, CONV2_RELU_F3out0 , LastRamOutF3_8 );
OneRegisterOut RAMFilter3Combined9  (clk, Stage2_xwrite_5, CONV2_RELU_F3out1 , LastRamOutF3_9 );

OneRegisterOut RAMFilter3Combined10  (clk, Stage2_xwrite_1, CONV2_RELU_F3out10 , LastRamOutF3_10 );
OneRegisterOut RAMFilter3Combined11  (clk, Stage2_xwrite_1, CONV2_RELU_F3out11 , LastRamOutF3_11 );
OneRegisterOut RAMFilter3Combined12  (clk, Stage2_xwrite_2, CONV2_RELU_F3out10 , LastRamOutF3_12 );
OneRegisterOut RAMFilter3Combined13  (clk, Stage2_xwrite_2, CONV2_RELU_F3out11 , LastRamOutF3_13 );
OneRegisterOut RAMFilter3Combined14  (clk, Stage2_xwrite_3, CONV2_RELU_F3out10 , LastRamOutF3_14 );
OneRegisterOut RAMFilter3Combined15  (clk, Stage2_xwrite_3, CONV2_RELU_F3out11 , LastRamOutF3_15 );
OneRegisterOut RAMFilter3Combined16  (clk, Stage2_xwrite_4, CONV2_RELU_F3out10 , LastRamOutF3_16 );
OneRegisterOut RAMFilter3Combined17  (clk, Stage2_xwrite_4, CONV2_RELU_F3out11 , LastRamOutF3_17 );
OneRegisterOut RAMFilter3Combined18  (clk, Stage2_xwrite_5, CONV2_RELU_F3out10 , LastRamOutF3_18 );
OneRegisterOut RAMFilter3Combined19  (clk, Stage2_xwrite_5, CONV2_RELU_F3out11 , LastRamOutF3_19 );

OneRegisterOut RAMFilter3Combined20  (clk, Stage2_xwrite_6, CONV2_RELU_F3out0 , LastRamOutF3_20 );
OneRegisterOut RAMFilter3Combined21  (clk, Stage2_xwrite_6, CONV2_RELU_F3out1 , LastRamOutF3_21 );
OneRegisterOut RAMFilter3Combined22  (clk, Stage2_xwrite_7, CONV2_RELU_F3out0 , LastRamOutF3_22 );
OneRegisterOut RAMFilter3Combined23  (clk, Stage2_xwrite_7, CONV2_RELU_F3out1 , LastRamOutF3_23 );
OneRegisterOut RAMFilter3Combined24  (clk, Stage2_xwrite_8, CONV2_RELU_F3out0 , LastRamOutF3_24 );
OneRegisterOut RAMFilter3Combined25  (clk, Stage2_xwrite_8, CONV2_RELU_F3out1 , LastRamOutF3_25 );
OneRegisterOut RAMFilter3Combined26  (clk, Stage2_xwrite_9, CONV2_RELU_F3out0 , LastRamOutF3_26 );
OneRegisterOut RAMFilter3Combined27  (clk, Stage2_xwrite_9, CONV2_RELU_F3out1 , LastRamOutF3_27 );
OneRegisterOut RAMFilter3Combined28  (clk, Stage2_xwrite_10, CONV2_RELU_F3out0 , LastRamOutF3_28 );
OneRegisterOut RAMFilter3Combined29  (clk, Stage2_xwrite_10, CONV2_RELU_F3out1 , LastRamOutF3_29 );

OneRegisterOut RAMFilter3Combined30  (clk, Stage2_xwrite_6, CONV2_RELU_F3out10 , LastRamOutF3_30 );
OneRegisterOut RAMFilter3Combined31  (clk, Stage2_xwrite_6, CONV2_RELU_F3out11 , LastRamOutF3_31 );
OneRegisterOut RAMFilter3Combined32  (clk, Stage2_xwrite_7, CONV2_RELU_F3out10 , LastRamOutF3_32 );
OneRegisterOut RAMFilter3Combined33  (clk, Stage2_xwrite_7, CONV2_RELU_F3out11 , LastRamOutF3_33 );
OneRegisterOut RAMFilter3Combined34  (clk, Stage2_xwrite_8, CONV2_RELU_F3out10 , LastRamOutF3_34 );
OneRegisterOut RAMFilter3Combined35  (clk, Stage2_xwrite_8, CONV2_RELU_F3out11 , LastRamOutF3_35 );
OneRegisterOut RAMFilter3Combined36  (clk, Stage2_xwrite_9, CONV2_RELU_F3out10 , LastRamOutF3_36 );
OneRegisterOut RAMFilter3Combined37  (clk, Stage2_xwrite_9, CONV2_RELU_F3out11 , LastRamOutF3_37 );
OneRegisterOut RAMFilter3Combined38  (clk, Stage2_xwrite_10, CONV2_RELU_F3out10 , LastRamOutF3_38 );
OneRegisterOut RAMFilter3Combined39  (clk, Stage2_xwrite_10, CONV2_RELU_F3out11 , LastRamOutF3_39 );

OneRegisterOut RAMFilter3Combined40  (clk, Stage2_xwrite_11, CONV2_RELU_F3out0 , LastRamOutF3_40 );
OneRegisterOut RAMFilter3Combined41  (clk, Stage2_xwrite_11, CONV2_RELU_F3out1 , LastRamOutF3_41 );
OneRegisterOut RAMFilter3Combined42  (clk, Stage2_xwrite_12, CONV2_RELU_F3out0 , LastRamOutF3_42 );
OneRegisterOut RAMFilter3Combined43  (clk, Stage2_xwrite_12, CONV2_RELU_F3out1 , LastRamOutF3_43 );
OneRegisterOut RAMFilter3Combined44  (clk, Stage2_xwrite_13, CONV2_RELU_F3out0 , LastRamOutF3_44 );
OneRegisterOut RAMFilter3Combined45  (clk, Stage2_xwrite_13, CONV2_RELU_F3out1 , LastRamOutF3_45 );
OneRegisterOut RAMFilter3Combined46  (clk, Stage2_xwrite_14, CONV2_RELU_F3out0 , LastRamOutF3_46 );
OneRegisterOut RAMFilter3Combined47  (clk, Stage2_xwrite_14, CONV2_RELU_F3out1 , LastRamOutF3_47 );
OneRegisterOut RAMFilter3Combined48  (clk, Stage2_xwrite_15, CONV2_RELU_F3out0 , LastRamOutF3_48 );
OneRegisterOut RAMFilter3Combined49  (clk, Stage2_xwrite_15, CONV2_RELU_F3out1 , LastRamOutF3_49 );

OneRegisterOut RAMFilter3Combined50  (clk, Stage2_xwrite_11, CONV2_RELU_F3out10 , LastRamOutF3_50 );
OneRegisterOut RAMFilter3Combined51  (clk, Stage2_xwrite_11, CONV2_RELU_F3out11 , LastRamOutF3_51 );
OneRegisterOut RAMFilter3Combined52  (clk, Stage2_xwrite_12, CONV2_RELU_F3out10 , LastRamOutF3_52 );
OneRegisterOut RAMFilter3Combined53  (clk, Stage2_xwrite_12, CONV2_RELU_F3out11 , LastRamOutF3_53 );
OneRegisterOut RAMFilter3Combined54  (clk, Stage2_xwrite_13, CONV2_RELU_F3out10 , LastRamOutF3_54 );
OneRegisterOut RAMFilter3Combined55  (clk, Stage2_xwrite_13, CONV2_RELU_F3out11 , LastRamOutF3_55 );
OneRegisterOut RAMFilter3Combined56  (clk, Stage2_xwrite_14, CONV2_RELU_F3out10 , LastRamOutF3_56 );
OneRegisterOut RAMFilter3Combined57  (clk, Stage2_xwrite_14, CONV2_RELU_F3out11 , LastRamOutF3_57 );
OneRegisterOut RAMFilter3Combined58  (clk, Stage2_xwrite_15, CONV2_RELU_F3out10 , LastRamOutF3_58 );
OneRegisterOut RAMFilter3Combined59  (clk, Stage2_xwrite_15, CONV2_RELU_F3out11 , LastRamOutF3_59 );

OneRegisterOut RAMFilter3Combined60  (clk, Stage2_xwrite_16, CONV2_RELU_F3out0 , LastRamOutF3_60 );
OneRegisterOut RAMFilter3Combined61  (clk, Stage2_xwrite_16, CONV2_RELU_F3out1 , LastRamOutF3_61 );
OneRegisterOut RAMFilter3Combined62  (clk, Stage2_xwrite_17, CONV2_RELU_F3out0 , LastRamOutF3_62 );
OneRegisterOut RAMFilter3Combined63  (clk, Stage2_xwrite_17, CONV2_RELU_F3out1 , LastRamOutF3_63 );
OneRegisterOut RAMFilter3Combined64  (clk, Stage2_xwrite_18, CONV2_RELU_F3out0 , LastRamOutF3_64 );
OneRegisterOut RAMFilter3Combined65  (clk, Stage2_xwrite_18, CONV2_RELU_F3out1 , LastRamOutF3_65 );
OneRegisterOut RAMFilter3Combined66  (clk, Stage2_xwrite_19, CONV2_RELU_F3out0 , LastRamOutF3_66 );
OneRegisterOut RAMFilter3Combined67  (clk, Stage2_xwrite_19, CONV2_RELU_F3out1 , LastRamOutF3_67 );
OneRegisterOut RAMFilter3Combined68  (clk, Stage2_xwrite_20, CONV2_RELU_F3out0 , LastRamOutF3_68 );
OneRegisterOut RAMFilter3Combined69  (clk, Stage2_xwrite_20, CONV2_RELU_F3out1 , LastRamOutF3_69 );

OneRegisterOut RAMFilter3Combined70  (clk, Stage2_xwrite_16, CONV2_RELU_F3out10 , LastRamOutF3_70 );
OneRegisterOut RAMFilter3Combined71  (clk, Stage2_xwrite_16, CONV2_RELU_F3out11 , LastRamOutF3_71 );
OneRegisterOut RAMFilter3Combined72  (clk, Stage2_xwrite_17, CONV2_RELU_F3out10 , LastRamOutF3_72 );
OneRegisterOut RAMFilter3Combined73  (clk, Stage2_xwrite_17, CONV2_RELU_F3out11 , LastRamOutF3_73 );
OneRegisterOut RAMFilter3Combined74  (clk, Stage2_xwrite_18, CONV2_RELU_F3out10 , LastRamOutF3_74 );
OneRegisterOut RAMFilter3Combined75  (clk, Stage2_xwrite_18, CONV2_RELU_F3out11 , LastRamOutF3_75 );
OneRegisterOut RAMFilter3Combined76  (clk, Stage2_xwrite_19, CONV2_RELU_F3out10 , LastRamOutF3_76 );
OneRegisterOut RAMFilter3Combined77  (clk, Stage2_xwrite_19, CONV2_RELU_F3out11 , LastRamOutF3_77 );
OneRegisterOut RAMFilter3Combined78  (clk, Stage2_xwrite_20, CONV2_RELU_F3out10 , LastRamOutF3_78 );
OneRegisterOut RAMFilter3Combined79  (clk, Stage2_xwrite_20, CONV2_RELU_F3out11 , LastRamOutF3_79 );

OneRegisterOut RAMFilter3Combined80  (clk, Stage2_xwrite_21, CONV2_RELU_F3out0 , LastRamOutF3_80 );
OneRegisterOut RAMFilter3Combined81  (clk, Stage2_xwrite_21, CONV2_RELU_F3out1 , LastRamOutF3_81 );
OneRegisterOut RAMFilter3Combined82  (clk, Stage2_xwrite_22, CONV2_RELU_F3out0 , LastRamOutF3_82 );
OneRegisterOut RAMFilter3Combined83  (clk, Stage2_xwrite_22, CONV2_RELU_F3out1 , LastRamOutF3_83 );
OneRegisterOut RAMFilter3Combined84  (clk, Stage2_xwrite_23, CONV2_RELU_F3out0 , LastRamOutF3_84 );
OneRegisterOut RAMFilter3Combined85  (clk, Stage2_xwrite_23, CONV2_RELU_F3out1 , LastRamOutF3_85 );
OneRegisterOut RAMFilter3Combined86  (clk, Stage2_xwrite_24, CONV2_RELU_F3out0 , LastRamOutF3_86 );
OneRegisterOut RAMFilter3Combined87  (clk, Stage2_xwrite_24, CONV2_RELU_F3out1 , LastRamOutF3_87 );
OneRegisterOut RAMFilter3Combined88  (clk, Stage2_xwrite_25, CONV2_RELU_F3out0 , LastRamOutF3_88 );
OneRegisterOut RAMFilter3Combined89  (clk, Stage2_xwrite_25, CONV2_RELU_F3out1 , LastRamOutF3_89 );

OneRegisterOut RAMFilter3Combined90  (clk, Stage2_xwrite_21, CONV2_RELU_F3out10 , LastRamOutF3_90 );
OneRegisterOut RAMFilter3Combined91  (clk, Stage2_xwrite_21, CONV2_RELU_F3out11 , LastRamOutF3_91 );
OneRegisterOut RAMFilter3Combined92  (clk, Stage2_xwrite_22, CONV2_RELU_F3out10 , LastRamOutF3_92 );
OneRegisterOut RAMFilter3Combined93  (clk, Stage2_xwrite_22, CONV2_RELU_F3out11 , LastRamOutF3_93 );
OneRegisterOut RAMFilter3Combined94  (clk, Stage2_xwrite_23, CONV2_RELU_F3out10 , LastRamOutF3_94 );
OneRegisterOut RAMFilter3Combined95  (clk, Stage2_xwrite_23, CONV2_RELU_F3out11 , LastRamOutF3_95 );
OneRegisterOut RAMFilter3Combined96  (clk, Stage2_xwrite_24, CONV2_RELU_F3out10 , LastRamOutF3_96 );
OneRegisterOut RAMFilter3Combined97  (clk, Stage2_xwrite_24, CONV2_RELU_F3out11 , LastRamOutF3_97 );
OneRegisterOut RAMFilter3Combined98  (clk, Stage2_xwrite_25, CONV2_RELU_F3out10 , LastRamOutF3_98 );
OneRegisterOut RAMFilter3Combined99  (clk, Stage2_xwrite_25, CONV2_RELU_F3out11 , LastRamOutF3_99 );

////



OneRegisterOut RAMFilter4Combined0  (clk, Stage2_xwrite_1, CONV2_RELU_F4out0 , LastRamOutF4_0 );
OneRegisterOut RAMFilter4Combined1  (clk, Stage2_xwrite_1, CONV2_RELU_F4out1 , LastRamOutF4_1 );
OneRegisterOut RAMFilter4Combined2  (clk, Stage2_xwrite_2, CONV2_RELU_F4out0 , LastRamOutF4_2 );
OneRegisterOut RAMFilter4Combined3  (clk, Stage2_xwrite_2, CONV2_RELU_F4out1 , LastRamOutF4_3 );
OneRegisterOut RAMFilter4Combined4  (clk, Stage2_xwrite_3, CONV2_RELU_F4out0 , LastRamOutF4_4 );
OneRegisterOut RAMFilter4Combined5  (clk, Stage2_xwrite_3, CONV2_RELU_F4out1 , LastRamOutF4_5 );
OneRegisterOut RAMFilter4Combined6  (clk, Stage2_xwrite_4, CONV2_RELU_F4out0 , LastRamOutF4_6 );
OneRegisterOut RAMFilter4Combined7  (clk, Stage2_xwrite_4, CONV2_RELU_F4out1 , LastRamOutF4_7 );
OneRegisterOut RAMFilter4Combined8  (clk, Stage2_xwrite_5, CONV2_RELU_F4out0 , LastRamOutF4_8 );
OneRegisterOut RAMFilter4Combined9  (clk, Stage2_xwrite_5, CONV2_RELU_F4out1 , LastRamOutF4_9 );

OneRegisterOut RAMFilter4Combined10  (clk, Stage2_xwrite_1, CONV2_RELU_F4out10 , LastRamOutF4_10 );
OneRegisterOut RAMFilter4Combined11  (clk, Stage2_xwrite_1, CONV2_RELU_F4out11 , LastRamOutF4_11 );
OneRegisterOut RAMFilter4Combined12  (clk, Stage2_xwrite_2, CONV2_RELU_F4out10 , LastRamOutF4_12 );
OneRegisterOut RAMFilter4Combined13  (clk, Stage2_xwrite_2, CONV2_RELU_F4out11 , LastRamOutF4_13 );
OneRegisterOut RAMFilter4Combined14  (clk, Stage2_xwrite_3, CONV2_RELU_F4out10 , LastRamOutF4_14 );
OneRegisterOut RAMFilter4Combined15  (clk, Stage2_xwrite_3, CONV2_RELU_F4out11 , LastRamOutF4_15 );
OneRegisterOut RAMFilter4Combined16  (clk, Stage2_xwrite_4, CONV2_RELU_F4out10 , LastRamOutF4_16 );
OneRegisterOut RAMFilter4Combined17  (clk, Stage2_xwrite_4, CONV2_RELU_F4out11 , LastRamOutF4_17 );
OneRegisterOut RAMFilter4Combined18  (clk, Stage2_xwrite_5, CONV2_RELU_F4out10 , LastRamOutF4_18 );
OneRegisterOut RAMFilter4Combined19  (clk, Stage2_xwrite_5, CONV2_RELU_F4out11 , LastRamOutF4_19 );

OneRegisterOut RAMFilter4Combined20  (clk, Stage2_xwrite_6, CONV2_RELU_F4out0 , LastRamOutF4_20 );
OneRegisterOut RAMFilter4Combined21  (clk, Stage2_xwrite_6, CONV2_RELU_F4out1 , LastRamOutF4_21 );
OneRegisterOut RAMFilter4Combined22  (clk, Stage2_xwrite_7, CONV2_RELU_F4out0 , LastRamOutF4_22 );
OneRegisterOut RAMFilter4Combined23  (clk, Stage2_xwrite_7, CONV2_RELU_F4out1 , LastRamOutF4_23 );
OneRegisterOut RAMFilter4Combined24  (clk, Stage2_xwrite_8, CONV2_RELU_F4out0 , LastRamOutF4_24 );
OneRegisterOut RAMFilter4Combined25  (clk, Stage2_xwrite_8, CONV2_RELU_F4out1 , LastRamOutF4_25 );
OneRegisterOut RAMFilter4Combined26  (clk, Stage2_xwrite_9, CONV2_RELU_F4out0 , LastRamOutF4_26 );
OneRegisterOut RAMFilter4Combined27  (clk, Stage2_xwrite_9, CONV2_RELU_F4out1 , LastRamOutF4_27 );
OneRegisterOut RAMFilter4Combined28  (clk, Stage2_xwrite_10, CONV2_RELU_F4out0 , LastRamOutF4_28 );
OneRegisterOut RAMFilter4Combined29  (clk, Stage2_xwrite_10, CONV2_RELU_F4out1 , LastRamOutF4_29 );

OneRegisterOut RAMFilter4Combined30  (clk, Stage2_xwrite_6, CONV2_RELU_F4out10 , LastRamOutF4_30 );
OneRegisterOut RAMFilter4Combined31  (clk, Stage2_xwrite_6, CONV2_RELU_F4out11 , LastRamOutF4_31 );
OneRegisterOut RAMFilter4Combined32  (clk, Stage2_xwrite_7, CONV2_RELU_F4out10 , LastRamOutF4_32 );
OneRegisterOut RAMFilter4Combined33  (clk, Stage2_xwrite_7, CONV2_RELU_F4out11 , LastRamOutF4_33 );
OneRegisterOut RAMFilter4Combined34  (clk, Stage2_xwrite_8, CONV2_RELU_F4out10 , LastRamOutF4_34 );
OneRegisterOut RAMFilter4Combined35  (clk, Stage2_xwrite_8, CONV2_RELU_F4out11 , LastRamOutF4_35 );
OneRegisterOut RAMFilter4Combined36  (clk, Stage2_xwrite_9, CONV2_RELU_F4out10 , LastRamOutF4_36 );
OneRegisterOut RAMFilter4Combined37  (clk, Stage2_xwrite_9, CONV2_RELU_F4out11 , LastRamOutF4_37 );
OneRegisterOut RAMFilter4Combined38  (clk, Stage2_xwrite_10, CONV2_RELU_F4out10 , LastRamOutF4_38 );
OneRegisterOut RAMFilter4Combined39  (clk, Stage2_xwrite_10, CONV2_RELU_F4out11 , LastRamOutF4_39 );

OneRegisterOut RAMFilter4Combined40  (clk, Stage2_xwrite_11, CONV2_RELU_F4out0 , LastRamOutF4_40 );
OneRegisterOut RAMFilter4Combined41  (clk, Stage2_xwrite_11, CONV2_RELU_F4out1 , LastRamOutF4_41 );
OneRegisterOut RAMFilter4Combined42  (clk, Stage2_xwrite_12, CONV2_RELU_F4out0 , LastRamOutF4_42 );
OneRegisterOut RAMFilter4Combined43  (clk, Stage2_xwrite_12, CONV2_RELU_F4out1 , LastRamOutF4_43 );
OneRegisterOut RAMFilter4Combined44  (clk, Stage2_xwrite_13, CONV2_RELU_F4out0 , LastRamOutF4_44 );
OneRegisterOut RAMFilter4Combined45  (clk, Stage2_xwrite_13, CONV2_RELU_F4out1 , LastRamOutF4_45 );
OneRegisterOut RAMFilter4Combined46  (clk, Stage2_xwrite_14, CONV2_RELU_F4out0 , LastRamOutF4_46 );
OneRegisterOut RAMFilter4Combined47  (clk, Stage2_xwrite_14, CONV2_RELU_F4out1 , LastRamOutF4_47 );
OneRegisterOut RAMFilter4Combined48  (clk, Stage2_xwrite_15, CONV2_RELU_F4out0 , LastRamOutF4_48 );
OneRegisterOut RAMFilter4Combined49  (clk, Stage2_xwrite_15, CONV2_RELU_F4out1 , LastRamOutF4_49 );

OneRegisterOut RAMFilter4Combined50  (clk, Stage2_xwrite_11, CONV2_RELU_F4out10 , LastRamOutF4_50 );
OneRegisterOut RAMFilter4Combined51  (clk, Stage2_xwrite_11, CONV2_RELU_F4out11 , LastRamOutF4_51 );
OneRegisterOut RAMFilter4Combined52  (clk, Stage2_xwrite_12, CONV2_RELU_F4out10 , LastRamOutF4_52 );
OneRegisterOut RAMFilter4Combined53  (clk, Stage2_xwrite_12, CONV2_RELU_F4out11 , LastRamOutF4_53 );
OneRegisterOut RAMFilter4Combined54  (clk, Stage2_xwrite_13, CONV2_RELU_F4out10 , LastRamOutF4_54 );
OneRegisterOut RAMFilter4Combined55  (clk, Stage2_xwrite_13, CONV2_RELU_F4out11 , LastRamOutF4_55 );
OneRegisterOut RAMFilter4Combined56  (clk, Stage2_xwrite_14, CONV2_RELU_F4out10 , LastRamOutF4_56 );
OneRegisterOut RAMFilter4Combined57  (clk, Stage2_xwrite_14, CONV2_RELU_F4out11 , LastRamOutF4_57 );
OneRegisterOut RAMFilter4Combined58  (clk, Stage2_xwrite_15, CONV2_RELU_F4out10 , LastRamOutF4_58 );
OneRegisterOut RAMFilter4Combined59  (clk, Stage2_xwrite_15, CONV2_RELU_F4out11 , LastRamOutF4_59 );

OneRegisterOut RAMFilter4Combined60  (clk, Stage2_xwrite_16, CONV2_RELU_F4out0 , LastRamOutF4_60 );
OneRegisterOut RAMFilter4Combined61  (clk, Stage2_xwrite_16, CONV2_RELU_F4out1 , LastRamOutF4_61 );
OneRegisterOut RAMFilter4Combined62  (clk, Stage2_xwrite_17, CONV2_RELU_F4out0 , LastRamOutF4_62 );
OneRegisterOut RAMFilter4Combined63  (clk, Stage2_xwrite_17, CONV2_RELU_F4out1 , LastRamOutF4_63 );
OneRegisterOut RAMFilter4Combined64  (clk, Stage2_xwrite_18, CONV2_RELU_F4out0 , LastRamOutF4_64 );
OneRegisterOut RAMFilter4Combined65  (clk, Stage2_xwrite_18, CONV2_RELU_F4out1 , LastRamOutF4_65 );
OneRegisterOut RAMFilter4Combined66  (clk, Stage2_xwrite_19, CONV2_RELU_F4out0 , LastRamOutF4_66 );
OneRegisterOut RAMFilter4Combined67  (clk, Stage2_xwrite_19, CONV2_RELU_F4out1 , LastRamOutF4_67 );
OneRegisterOut RAMFilter4Combined68  (clk, Stage2_xwrite_20, CONV2_RELU_F4out0 , LastRamOutF4_68 );
OneRegisterOut RAMFilter4Combined69  (clk, Stage2_xwrite_20, CONV2_RELU_F4out1 , LastRamOutF4_69 );

OneRegisterOut RAMFilter4Combined70  (clk, Stage2_xwrite_16, CONV2_RELU_F4out10 , LastRamOutF4_70 );
OneRegisterOut RAMFilter4Combined71  (clk, Stage2_xwrite_16, CONV2_RELU_F4out11 , LastRamOutF4_71 );
OneRegisterOut RAMFilter4Combined72  (clk, Stage2_xwrite_17, CONV2_RELU_F4out10 , LastRamOutF4_72 );
OneRegisterOut RAMFilter4Combined73  (clk, Stage2_xwrite_17, CONV2_RELU_F4out11 , LastRamOutF4_73 );
OneRegisterOut RAMFilter4Combined74  (clk, Stage2_xwrite_18, CONV2_RELU_F4out10 , LastRamOutF4_74 );
OneRegisterOut RAMFilter4Combined75  (clk, Stage2_xwrite_18, CONV2_RELU_F4out11 , LastRamOutF4_75 );
OneRegisterOut RAMFilter4Combined76  (clk, Stage2_xwrite_19, CONV2_RELU_F4out10 , LastRamOutF4_76 );
OneRegisterOut RAMFilter4Combined77  (clk, Stage2_xwrite_19, CONV2_RELU_F4out11 , LastRamOutF4_77 );
OneRegisterOut RAMFilter4Combined78  (clk, Stage2_xwrite_20, CONV2_RELU_F4out10 , LastRamOutF4_78 );
OneRegisterOut RAMFilter4Combined79  (clk, Stage2_xwrite_20, CONV2_RELU_F4out11 , LastRamOutF4_79 );

OneRegisterOut RAMFilter4Combined80  (clk, Stage2_xwrite_21, CONV2_RELU_F4out0 , LastRamOutF4_80 );
OneRegisterOut RAMFilter4Combined81  (clk, Stage2_xwrite_21, CONV2_RELU_F4out1 , LastRamOutF4_81 );
OneRegisterOut RAMFilter4Combined82  (clk, Stage2_xwrite_22, CONV2_RELU_F4out0 , LastRamOutF4_82 );
OneRegisterOut RAMFilter4Combined83  (clk, Stage2_xwrite_22, CONV2_RELU_F4out1 , LastRamOutF4_83 );
OneRegisterOut RAMFilter4Combined84  (clk, Stage2_xwrite_23, CONV2_RELU_F4out0 , LastRamOutF4_84 );
OneRegisterOut RAMFilter4Combined85  (clk, Stage2_xwrite_23, CONV2_RELU_F4out1 , LastRamOutF4_85 );
OneRegisterOut RAMFilter4Combined86  (clk, Stage2_xwrite_24, CONV2_RELU_F4out0 , LastRamOutF4_86 );
OneRegisterOut RAMFilter4Combined87  (clk, Stage2_xwrite_24, CONV2_RELU_F4out1 , LastRamOutF4_87 );
OneRegisterOut RAMFilter4Combined88  (clk, Stage2_xwrite_25, CONV2_RELU_F4out0 , LastRamOutF4_88 );
OneRegisterOut RAMFilter4Combined89  (clk, Stage2_xwrite_25, CONV2_RELU_F4out1 , LastRamOutF4_89 );

OneRegisterOut RAMFilter4Combined90  (clk, Stage2_xwrite_21, CONV2_RELU_F4out10 , LastRamOutF4_90 );
OneRegisterOut RAMFilter4Combined91  (clk, Stage2_xwrite_21, CONV2_RELU_F4out11 , LastRamOutF4_91 );
OneRegisterOut RAMFilter4Combined92  (clk, Stage2_xwrite_22, CONV2_RELU_F4out10 , LastRamOutF4_92 );
OneRegisterOut RAMFilter4Combined93  (clk, Stage2_xwrite_22, CONV2_RELU_F4out11 , LastRamOutF4_93 );
OneRegisterOut RAMFilter4Combined94  (clk, Stage2_xwrite_23, CONV2_RELU_F4out10 , LastRamOutF4_94 );
OneRegisterOut RAMFilter4Combined95  (clk, Stage2_xwrite_23, CONV2_RELU_F4out11 , LastRamOutF4_95 );
OneRegisterOut RAMFilter4Combined96  (clk, Stage2_xwrite_24, CONV2_RELU_F4out10 , LastRamOutF4_96 );
OneRegisterOut RAMFilter4Combined97  (clk, Stage2_xwrite_24, CONV2_RELU_F4out11 , LastRamOutF4_97 );
OneRegisterOut RAMFilter4Combined98  (clk, Stage2_xwrite_25, CONV2_RELU_F4out10 , LastRamOutF4_98 );
OneRegisterOut RAMFilter4Combined99  (clk, Stage2_xwrite_25, CONV2_RELU_F4out11 , LastRamOutF4_99 );

endmodule
*/