module TB_bla();

reg clk;
reg rst_Controller;
//reg L0START;
//wire L0FINISH;
reg [65:0] DataIn0 , DataIn1 , DataIn2 , DataIn3 ;

localparam period = 100; 
/* wire [65:0] FinalAnswer; */
wire [3:0] FinalAnswer;
//LAYER0 TheLayer(clk ,L0START, L0FINISH , DataIn0 , DataIn1 , DataIn2 , DataIn3 , DataOut0 , DataOut1 , DataOut2 , DataOut3 , DataOut4 , DataOut5 , DataOut6 , DataOut7 , DataOut8 , DataOut9 , DataOut10 , DataOut11 , DataOut12 , DataOut13 , DataOut14 , DataOut15 , DataOut16 , DataOut17 , DataOut18 , DataOut19 , DataOut20 , DataOut21 , DataOut22 , DataOut23 , DataOut24 , DataOut25 , DataOut26 , DataOut27 , DataOut28 , DataOut29 , DataOut30 , DataOut31 , DataOut32 , DataOut33 , DataOut34 , DataOut35 , DataOut36 , DataOut37 , DataOut38 , DataOut39 , DataOut40 , DataOut41 , DataOut42 , DataOut43 , DataOut44 , DataOut45 , DataOut46 , DataOut47 , DataOut48 , DataOut49 , DataOut50 , DataOut51 , DataOut52 , DataOut53 , DataOut54 , DataOut55 , DataOut56 , DataOut57 , DataOut58 , DataOut59 , DataOut60 , DataOut61 , DataOut62 , DataOut63 , DataOut64 , DataOut65 , DataOut66 , DataOut67 , DataOut68 , DataOut69 , DataOut70 , DataOut71 , DataOut72 , DataOut73 , DataOut74 , DataOut75 , DataOut76 , DataOut77 , DataOut78 , DataOut79 , DataOut80 , DataOut81 , DataOut82 , DataOut83 , DataOut84 , DataOut85 , DataOut86 , DataOut87 , DataOut88 , DataOut89 , DataOut90 , DataOut91 , DataOut92 , DataOut93 , DataOut94 , DataOut95 , DataOut96 , DataOut97 , DataOut98 , DataOut99 , DataOut100 , DataOut101 , DataOut102 , DataOut103 , DataOut104 , DataOut105 , DataOut106 , DataOut107 , DataOut108 , DataOut109 , DataOut110 , DataOut111 , DataOut112 , DataOut113 , DataOut114 , DataOut115 , DataOut116 , DataOut117 , DataOut118 , DataOut119 , DataOut120 , DataOut121 , DataOut122 , DataOut123 , DataOut124 , DataOut125 , DataOut126 , DataOut127 , DataOut128 , DataOut129 , DataOut130 , DataOut131 , DataOut132 , DataOut133 , DataOut134 , DataOut135 , DataOut136 , DataOut137 , DataOut138 , DataOut139 , DataOut140 , DataOut141 , DataOut142 , DataOut143 , DataOut144 , DataOut145 , DataOut146 , DataOut147 , DataOut148 , DataOut149 , DataOut150 , DataOut151 , DataOut152 , DataOut153 , DataOut154 , DataOut155 , DataOut156 , DataOut157 , DataOut158 , DataOut159 , DataOut160 , DataOut161 , DataOut162 , DataOut163 , DataOut164 , DataOut165 , DataOut166 , DataOut167 , DataOut168 , DataOut169 , DataOut170 , DataOut171 , DataOut172 , DataOut173 , DataOut174 , DataOut175 , DataOut176 , DataOut177 , DataOut178 , DataOut179 , DataOut180 , DataOut181 , DataOut182 , DataOut183 , DataOut184 , DataOut185 , DataOut186 , DataOut187 , DataOut188 , DataOut189 , DataOut190 , DataOut191 , DataOut192 , DataOut193 , DataOut194 , DataOut195 , DataOut196 , DataOut197 , DataOut198 , DataOut199 , DataOut200 , DataOut201 , DataOut202 , DataOut203 , DataOut204 , DataOut205 , DataOut206 , DataOut207 , DataOut208 , DataOut209 , DataOut210 , DataOut211 , DataOut212 , DataOut213 , DataOut214 , DataOut215 , DataOut216 , DataOut217 , DataOut218 , DataOut219 , DataOut220 , DataOut221 , DataOut222 , DataOut223 , DataOut224 , DataOut225 , DataOut226 , DataOut227 , DataOut228 , DataOut229 , DataOut230 , DataOut231 , DataOut232 , DataOut233 , DataOut234 , DataOut235 , DataOut236 , DataOut237 , DataOut238 , DataOut239 , DataOut240 , DataOut241 , DataOut242 , DataOut243 , DataOut244 , DataOut245 , DataOut246 , DataOut247 , DataOut248 , DataOut249 , DataOut250 , DataOut251 , DataOut252 , DataOut253 , DataOut254 , DataOut255 , DataOut256 , DataOut257 , DataOut258 , DataOut259 , DataOut260 , DataOut261 , DataOut262 , DataOut263 , DataOut264 , DataOut265 , DataOut266 , DataOut267 , DataOut268 , DataOut269 , DataOut270 , DataOut271 , DataOut272 , DataOut273 , DataOut274 , DataOut275 , DataOut276 , DataOut277 , DataOut278 , DataOut279 , DataOut280 , DataOut281 , DataOut282 , DataOut283 , DataOut284 , DataOut285 , DataOut286 , DataOut287 , DataOut288 , DataOut289 , DataOut290 , DataOut291 , DataOut292 , DataOut293 , DataOut294 , DataOut295 , DataOut296 , DataOut297 , DataOut298 , DataOut299 , DataOut300 , DataOut301 , DataOut302 , DataOut303 , DataOut304 , DataOut305 , DataOut306 , DataOut307 , DataOut308 , DataOut309 , DataOut310 , DataOut311 , DataOut312 , DataOut313 , DataOut314 , DataOut315 , DataOut316 , DataOut317 , DataOut318 , DataOut319 , DataOut320 , DataOut321 , DataOut322 , DataOut323 , DataOut324 , DataOut325 , DataOut326 , DataOut327 , DataOut328 , DataOut329 , DataOut330 , DataOut331 , DataOut332 , DataOut333 , DataOut334 , DataOut335 , DataOut336 , DataOut337 , DataOut338 , DataOut339 , DataOut340 , DataOut341 , DataOut342 , DataOut343 , DataOut344 , DataOut345 , DataOut346 , DataOut347 , DataOut348 , DataOut349 , DataOut350 , DataOut351 , DataOut352 , DataOut353 , DataOut354 , DataOut355 , DataOut356 , DataOut357 , DataOut358 , DataOut359 , DataOut360 , DataOut361 , DataOut362 , DataOut363 , DataOut364 , DataOut365 , DataOut366 , DataOut367 , DataOut368 , DataOut369 , DataOut370 , DataOut371 , DataOut372 , DataOut373 , DataOut374 , DataOut375 , DataOut376 , DataOut377 , DataOut378 , DataOut379 , DataOut380 , DataOut381 , DataOut382 , DataOut383 , DataOut384 , DataOut385 , DataOut386 , DataOut387 , DataOut388 , DataOut389 , DataOut390 , DataOut391 , DataOut392 , DataOut393 , DataOut394 , DataOut395 , DataOut396 , DataOut397 , DataOut398 , DataOut399 , DataOut400 , DataOut401 , DataOut402 , DataOut403 , DataOut404 , DataOut405 , DataOut406 , DataOut407 , DataOut408 , DataOut409 , DataOut410 , DataOut411 , DataOut412 , DataOut413 , DataOut414 , DataOut415 , DataOut416 , DataOut417 , DataOut418 , DataOut419 , DataOut420 , DataOut421 , DataOut422 , DataOut423 , DataOut424 , DataOut425 , DataOut426 , DataOut427 , DataOut428 , DataOut429 , DataOut430 , DataOut431 , DataOut432 , DataOut433 , DataOut434 , DataOut435 , DataOut436 , DataOut437 , DataOut438 , DataOut439 , DataOut440 , DataOut441 , DataOut442 , DataOut443 , DataOut444 , DataOut445 , DataOut446 , DataOut447 , DataOut448 , DataOut449 , DataOut450 , DataOut451 , DataOut452 , DataOut453 , DataOut454 , DataOut455 , DataOut456 , DataOut457 , DataOut458 , DataOut459 , DataOut460 , DataOut461 , DataOut462 , DataOut463 , DataOut464 , DataOut465 , DataOut466 , DataOut467 , DataOut468 , DataOut469 , DataOut470 , DataOut471 , DataOut472 , DataOut473 , DataOut474 , DataOut475 , DataOut476 , DataOut477 , DataOut478 , DataOut479 , DataOut480 , DataOut481 , DataOut482 , DataOut483 , DataOut484 , DataOut485 , DataOut486 , DataOut487 , DataOut488 , DataOut489 , DataOut490 , DataOut491 , DataOut492 , DataOut493 , DataOut494 , DataOut495 , DataOut496 , DataOut497 , DataOut498 , DataOut499 , DataOut500 , DataOut501 , DataOut502 , DataOut503 , DataOut504 , DataOut505 , DataOut506 , DataOut507 , DataOut508 , DataOut509 , DataOut510 , DataOut511 , DataOut512 , DataOut513 , DataOut514 , DataOut515 , DataOut516 , DataOut517 , DataOut518 , DataOut519 , DataOut520 , DataOut521 , DataOut522 , DataOut523 , DataOut524 , DataOut525 , DataOut526 , DataOut527 , DataOut528 , DataOut529 , DataOut530 , DataOut531 , DataOut532 , DataOut533 , DataOut534 , DataOut535 , DataOut536 , DataOut537 , DataOut538 , DataOut539 , DataOut540 , DataOut541 , DataOut542 , DataOut543 , DataOut544 , DataOut545 , DataOut546 , DataOut547 , DataOut548 , DataOut549 , DataOut550 , DataOut551 , DataOut552 , DataOut553 , DataOut554 , DataOut555 , DataOut556 , DataOut557 , DataOut558 , DataOut559 , DataOut560 , DataOut561 , DataOut562 , DataOut563 , DataOut564 , DataOut565 , DataOut566 , DataOut567 , DataOut568 , DataOut569 , DataOut570 , DataOut571 , DataOut572 , DataOut573 , DataOut574 , DataOut575 , DataOut576 , DataOut577 , DataOut578 , DataOut579 , DataOut580 , DataOut581 , DataOut582 , DataOut583 , DataOut584 , DataOut585 , DataOut586 , DataOut587 , DataOut588 , DataOut589 , DataOut590 , DataOut591 , DataOut592 , DataOut593 , DataOut594 , DataOut595 , DataOut596 , DataOut597 , DataOut598 , DataOut599 , DataOut600 , DataOut601 , DataOut602 , DataOut603 , DataOut604 , DataOut605 , DataOut606 , DataOut607 , DataOut608 , DataOut609 , DataOut610 , DataOut611 , DataOut612 , DataOut613 , DataOut614 , DataOut615 , DataOut616 , DataOut617 , DataOut618 , DataOut619 , DataOut620 , DataOut621 , DataOut622 , DataOut623 , DataOut624 , DataOut625 , DataOut626 , DataOut627 , DataOut628 , DataOut629 , DataOut630 , DataOut631 , DataOut632 , DataOut633 , DataOut634 , DataOut635 , DataOut636 , DataOut637 , DataOut638 , DataOut639 , DataOut640 , DataOut641 , DataOut642 , DataOut643 , DataOut644 , DataOut645 , DataOut646 , DataOut647 , DataOut648 , DataOut649 , DataOut650 , DataOut651 , DataOut652 , DataOut653 , DataOut654 , DataOut655 , DataOut656 , DataOut657 , DataOut658 , DataOut659 , DataOut660 , DataOut661 , DataOut662 , DataOut663 , DataOut664 , DataOut665 , DataOut666 , DataOut667 , DataOut668 , DataOut669 , DataOut670 , DataOut671 , DataOut672 , DataOut673 , DataOut674 , DataOut675 , DataOut676 , DataOut677 , DataOut678 , DataOut679 , DataOut680 , DataOut681 , DataOut682 , DataOut683 , DataOut684 , DataOut685 , DataOut686 , DataOut687 , DataOut688 , DataOut689 , DataOut690 , DataOut691 , DataOut692 , DataOut693 , DataOut694 , DataOut695 , DataOut696 , DataOut697 , DataOut698 , DataOut699 , DataOut700 , DataOut701 , DataOut702 , DataOut703 , DataOut704 , DataOut705 , DataOut706 , DataOut707 , DataOut708 , DataOut709 , DataOut710 , DataOut711 , DataOut712 , DataOut713 , DataOut714 , DataOut715 , DataOut716 , DataOut717 , DataOut718 , DataOut719 , DataOut720 , DataOut721 , DataOut722 , DataOut723 , DataOut724 , DataOut725 , DataOut726 , DataOut727 , DataOut728 , DataOut729 , DataOut730 , DataOut731 , DataOut732 , DataOut733 , DataOut734 , DataOut735 , DataOut736 , DataOut737 , DataOut738 , DataOut739 , DataOut740 , DataOut741 , DataOut742 , DataOut743 , DataOut744 , DataOut745 , DataOut746 , DataOut747 , DataOut748 , DataOut749 , DataOut750 , DataOut751 , DataOut752 , DataOut753 , DataOut754 , DataOut755 , DataOut756 , DataOut757 , DataOut758 , DataOut759 , DataOut760 , DataOut761 , DataOut762 , DataOut763 , DataOut764 , DataOut765 , DataOut766 , DataOut767 , DataOut768 , DataOut769 , DataOut770 , DataOut771 , DataOut772 , DataOut773 , DataOut774 , DataOut775 , DataOut776 , DataOut777 , DataOut778 , DataOut779 , DataOut780 , DataOut781 , DataOut782 , DataOut783 );
happy  otta (clk, rst_Controller,FinalAnswer,  DataIn0 , DataIn1 , DataIn2 , DataIn3);
always 
begin
    clk = 1'b0; 
    #50; 

    clk = 1'b1;
    #50; 
end

initial 
        begin
		
	    rst_Controller = 1;
		#20;
		rst_Controller = 0;
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
//repeat first input again			
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
///
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000110010000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000111110000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001100001001000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100001001000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010101100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001010010000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010011111111110000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000101010000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010101100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111010000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101011001000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101110110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100010111000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000110000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001100110011000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101100111000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001001011000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000101110000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010010000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001011010000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001001110100000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001100111111000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001011011010000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001010100110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101000111000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101110011000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010101010000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100101100000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101001010000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001100010011000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001100010011000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001000110100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000100110000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000111101000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101001000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100101011000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010011111111110000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100101110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010110010000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001010000110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111100000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101010100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001010011000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001000111100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000111101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001010100110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100011001000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010100000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101110000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000111000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000111001000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101110000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100011001000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001100111010000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000011100000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001100100110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101100000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000101000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000101100000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000111101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010010110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000110001000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000110010000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000111101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001001000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000110001000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100100011000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000111101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001001000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000000110001000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010111100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101001000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000101000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000110000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101010001000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100010110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010011111111110000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000101110000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101001110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101001010000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010000100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000110101000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001100100001000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101110101000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000111111000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001001110000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101010100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101000010000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001001000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001001000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001000001000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001000100100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001001000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101010001000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100101011000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010101100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101110011000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101101001000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101110011000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001010101100000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001011100100000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101101111000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001010101100000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000100110000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000000101010000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001100110110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101110011000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001010001100000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000100000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001010011000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001100010010000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000001101111111000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000001101111110000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b010100000001101111111000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b010100000001100010010000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b010100000000110011000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b010100000000101110000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 
DataIn0   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn1   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn2   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
DataIn3   <=66'b000000000000000000000000000000000000000000000000000000000000000000 ;
#period; 


        end

endmodule



module LAYER0_bla (clk ,L0START, L0FINISH , DataIn0 , DataIn1 , DataIn2 , DataIn3 , DataOut448 , DataOut449 , DataOut450 , DataOut451 , DataOut452 , DataOut453 , DataOut454 , DataOut455 , DataOut456 , DataOut457 , DataOut458 , DataOut459 , DataOut460 , DataOut461 , DataOut462 , DataOut463 , DataOut464 , DataOut465 , DataOut466 , DataOut467 , DataOut468 , DataOut469 , DataOut470 , DataOut471 , DataOut472 , DataOut473 , DataOut474 , DataOut475 , DataOut476 , DataOut477 , DataOut478 , DataOut479 , DataOut480 , DataOut481 , DataOut482 , DataOut483 , DataOut484 , DataOut485 , DataOut486 , DataOut487 , DataOut488 , DataOut489 , DataOut490 , DataOut491 , DataOut492 , DataOut493 , DataOut494 , DataOut495 , DataOut496 , DataOut497 , DataOut498 , DataOut499 , DataOut500 , DataOut501 , DataOut502 , DataOut503 , DataOut504 , DataOut505 , DataOut506 , DataOut507 , DataOut508 , DataOut509 , DataOut510 , DataOut511 , DataOut512 , DataOut513 , DataOut514 , DataOut515 , DataOut516 , DataOut517 , DataOut518 , DataOut519 , DataOut520 , DataOut521 , DataOut522 , DataOut523 , DataOut524 , DataOut525 , DataOut526 , DataOut527 , DataOut528 , DataOut529 , DataOut530 , DataOut531 , DataOut532 , DataOut533 , DataOut534 , DataOut535 , DataOut536 , DataOut537 , DataOut538 , DataOut539 , DataOut540 , DataOut541 , DataOut542 , DataOut543 , DataOut544 , DataOut545 , DataOut546 , DataOut547 , DataOut548 , DataOut549 , DataOut550 , DataOut551 , DataOut552 , DataOut553 , DataOut554 , DataOut555 , DataOut556 , DataOut557 , DataOut558 , DataOut559 , DataOut560 , DataOut561 , DataOut562 , DataOut563 , DataOut564 , DataOut565 , DataOut566 , DataOut567 , DataOut568 , DataOut569 , DataOut570 , DataOut571 , DataOut572 , DataOut573 , DataOut574 , DataOut575 , DataOut576 , DataOut577 , DataOut578 , DataOut579 , DataOut580 , DataOut581 , DataOut582 , DataOut583 , DataOut584 , DataOut585 , DataOut586 , DataOut587 , DataOut588 , DataOut589 , DataOut590 , DataOut591 , DataOut592 , DataOut593 , DataOut594 , DataOut595 , DataOut596 , DataOut597 , DataOut598 , DataOut599 , DataOut600 , DataOut601 , DataOut602 , DataOut603 , DataOut604 , DataOut605 , DataOut606 , DataOut607 , DataOut608 , DataOut609 , DataOut610 , DataOut611 , DataOut612 , DataOut613 , DataOut614 , DataOut615 , DataOut616 , DataOut617 , DataOut618 , DataOut619 , DataOut620 , DataOut621 , DataOut622 , DataOut623 , DataOut624 , DataOut625 , DataOut626 , DataOut627 , DataOut628 , DataOut629 , DataOut630 , DataOut631 , DataOut632 , DataOut633 , DataOut634 , DataOut635 , DataOut636 , DataOut637 , DataOut638 , DataOut639 , DataOut640 , DataOut641 , DataOut642 , DataOut643 , DataOut644 , DataOut645 , DataOut646 , DataOut647 , DataOut648 , DataOut649 , DataOut650 , DataOut651 , DataOut652 , DataOut653 , DataOut654 , DataOut655 , DataOut656 , DataOut657 , DataOut658 , DataOut659 , DataOut660 , DataOut661 , DataOut662 , DataOut663 , DataOut664 , DataOut665 , DataOut666 , DataOut667 , DataOut668 , DataOut669 , DataOut670 , DataOut671 , DataOut672 , DataOut673 , DataOut674 , DataOut675 , DataOut676 , DataOut677 , DataOut678 , DataOut679 , DataOut680 , DataOut681 , DataOut682 , DataOut683 , DataOut684 , DataOut685 , DataOut686 , DataOut687 , DataOut688 , DataOut689 , DataOut690 , DataOut691 , DataOut692 , DataOut693 , DataOut694 , DataOut695 , DataOut696 , DataOut697 , DataOut698 , DataOut699 , DataOut700 , DataOut701 , DataOut702 , DataOut703 , DataOut704 , DataOut705 , DataOut706 , DataOut707 , DataOut708 , DataOut709 , DataOut710 , DataOut711 , DataOut712 , DataOut713 , DataOut714 , DataOut715 , DataOut716 , DataOut717 , DataOut718 , DataOut719 , DataOut720 , DataOut721 , DataOut722 , DataOut723 , DataOut724 , DataOut725 , DataOut726 , DataOut727 , DataOut728 , DataOut729 , DataOut730 , DataOut731 , DataOut732 , DataOut733 , DataOut734 , DataOut735 , DataOut736 , DataOut737 , DataOut738 , DataOut739 , DataOut740 , DataOut741 , DataOut742 , DataOut743 , DataOut744 , DataOut745 , DataOut746 , DataOut747 , DataOut748 , DataOut749 , DataOut750 , DataOut751 , DataOut752 , DataOut753 , DataOut754 , DataOut755 , DataOut756 , DataOut757 , DataOut758 , DataOut759 , DataOut760 , DataOut761 , DataOut762 , DataOut763 , DataOut764 , DataOut765 , DataOut766 , DataOut767 , DataOut768 , DataOut769 , DataOut770 , DataOut771 , DataOut772 , DataOut773 , DataOut774 , DataOut775 , DataOut776 , DataOut777 , DataOut778 , DataOut779 , DataOut780 , DataOut781 , DataOut782 , DataOut783 );

input clk;
output reg [65:0] DataOut448 , DataOut449 , DataOut450 , DataOut451 , DataOut452 , DataOut453 , DataOut454 , DataOut455 , DataOut456 , DataOut457 , DataOut458 , DataOut459 , DataOut460 , DataOut461 , DataOut462 , DataOut463 , DataOut464 , DataOut465 , DataOut466 , DataOut467 , DataOut468 , DataOut469 , DataOut470 , DataOut471 , DataOut472 , DataOut473 , DataOut474 , DataOut475 , DataOut476 , DataOut477 , DataOut478 , DataOut479 , DataOut480 , DataOut481 , DataOut482 , DataOut483 , DataOut484 , DataOut485 , DataOut486 , DataOut487 , DataOut488 , DataOut489 , DataOut490 , DataOut491 , DataOut492 , DataOut493 , DataOut494 , DataOut495 , DataOut496 , DataOut497 , DataOut498 , DataOut499 , DataOut500 , DataOut501 , DataOut502 , DataOut503 , DataOut504 , DataOut505 , DataOut506 , DataOut507 , DataOut508 , DataOut509 , DataOut510 , DataOut511 , DataOut512 , DataOut513 , DataOut514 , DataOut515 , DataOut516 , DataOut517 , DataOut518 , DataOut519 , DataOut520 , DataOut521 , DataOut522 , DataOut523 , DataOut524 , DataOut525 , DataOut526 , DataOut527 , DataOut528 , DataOut529 , DataOut530 , DataOut531 , DataOut532 , DataOut533 , DataOut534 , DataOut535 , DataOut536 , DataOut537 , DataOut538 , DataOut539 , DataOut540 , DataOut541 , DataOut542 , DataOut543 , DataOut544 , DataOut545 , DataOut546 , DataOut547 , DataOut548 , DataOut549 , DataOut550 , DataOut551 , DataOut552 , DataOut553 , DataOut554 , DataOut555 , DataOut556 , DataOut557 , DataOut558 , DataOut559 , DataOut560 , DataOut561 , DataOut562 , DataOut563 , DataOut564 , DataOut565 , DataOut566 , DataOut567 , DataOut568 , DataOut569 , DataOut570 , DataOut571 , DataOut572 , DataOut573 , DataOut574 , DataOut575 , DataOut576 , DataOut577 , DataOut578 , DataOut579 , DataOut580 , DataOut581 , DataOut582 , DataOut583 , DataOut584 , DataOut585 , DataOut586 , DataOut587 , DataOut588 , DataOut589 , DataOut590 , DataOut591 , DataOut592 , DataOut593 , DataOut594 , DataOut595 , DataOut596 , DataOut597 , DataOut598 , DataOut599 , DataOut600 , DataOut601 , DataOut602 , DataOut603 , DataOut604 , DataOut605 , DataOut606 , DataOut607 , DataOut608 , DataOut609 , DataOut610 , DataOut611 , DataOut612 , DataOut613 , DataOut614 , DataOut615 , DataOut616 , DataOut617 , DataOut618 , DataOut619 , DataOut620 , DataOut621 , DataOut622 , DataOut623 , DataOut624 , DataOut625 , DataOut626 , DataOut627 , DataOut628 , DataOut629 , DataOut630 , DataOut631 , DataOut632 , DataOut633 , DataOut634 , DataOut635 , DataOut636 , DataOut637 , DataOut638 , DataOut639 , DataOut640 , DataOut641 , DataOut642 , DataOut643 , DataOut644 , DataOut645 , DataOut646 , DataOut647 , DataOut648 , DataOut649 , DataOut650 , DataOut651 , DataOut652 , DataOut653 , DataOut654 , DataOut655 , DataOut656 , DataOut657 , DataOut658 , DataOut659 , DataOut660 , DataOut661 , DataOut662 , DataOut663 , DataOut664 , DataOut665 , DataOut666 , DataOut667 , DataOut668 , DataOut669 , DataOut670 , DataOut671 , DataOut672 , DataOut673 , DataOut674 , DataOut675 , DataOut676 , DataOut677 , DataOut678 , DataOut679 , DataOut680 , DataOut681 , DataOut682 , DataOut683 , DataOut684 , DataOut685 , DataOut686 , DataOut687 , DataOut688 , DataOut689 , DataOut690 , DataOut691 , DataOut692 , DataOut693 , DataOut694 , DataOut695 , DataOut696 , DataOut697 , DataOut698 , DataOut699 , DataOut700 , DataOut701 , DataOut702 , DataOut703 , DataOut704 , DataOut705 , DataOut706 , DataOut707 , DataOut708 , DataOut709 , DataOut710 , DataOut711 , DataOut712 , DataOut713 , DataOut714 , DataOut715 , DataOut716 , DataOut717 , DataOut718 , DataOut719 , DataOut720 , DataOut721 , DataOut722 , DataOut723 , DataOut724 , DataOut725 , DataOut726 , DataOut727 , DataOut728 , DataOut729 , DataOut730 , DataOut731 , DataOut732 , DataOut733 , DataOut734 , DataOut735 , DataOut736 , DataOut737 , DataOut738 , DataOut739 , DataOut740 , DataOut741 , DataOut742 , DataOut743 , DataOut744 , DataOut745 , DataOut746 , DataOut747 , DataOut748 , DataOut749 , DataOut750 , DataOut751 , DataOut752 , DataOut753 , DataOut754 , DataOut755 , DataOut756 , DataOut757 , DataOut758 , DataOut759 , DataOut760 , DataOut761 , DataOut762 , DataOut763 , DataOut764 , DataOut765 , DataOut766 , DataOut767 , DataOut768 , DataOut769 , DataOut770 , DataOut771 , DataOut772 , DataOut773 , DataOut774 , DataOut775 , DataOut776 , DataOut777 , DataOut778 , DataOut779 , DataOut780 , DataOut781 , DataOut782 , DataOut783  ;
input L0START;
output reg L0FINISH;
input wire [65:0] DataIn0 , DataIn1 , DataIn2 , DataIn3 ;
wire [6:0] counter; 
wire dump; 
COUNTER_LAYER_128_cycles TheCounter (clk, counter, L0START,dump);
//counter 196 cycles : 8 bits
always @(posedge clk) 
begin 

//$monitor("counter = %b, L0START = %b, L0FINISH = %b , DataIn0= %b", counter , L0START, L0FINISH, DataIn0);

if (L0START)
begin
//$display("one");

case(counter)
0 : begin DataOut448  <=  DataIn0; DataOut449  <=  DataIn1; DataOut450  <=  DataIn2; DataOut451  <=  DataIn3; end
1  : begin DataOut452  <=  DataIn0; DataOut453  <=  DataIn1; DataOut454  <=  DataIn2; DataOut455  <=  DataIn3; end
2  : begin DataOut456  <=  DataIn0; DataOut457  <=  DataIn1; DataOut458  <=  DataIn2; DataOut459  <=  DataIn3; end
3  : begin DataOut460  <=  DataIn0; DataOut461  <=  DataIn1; DataOut462  <=  DataIn2; DataOut463  <=  DataIn3; end
4  : begin DataOut464  <=  DataIn0; DataOut465  <=  DataIn1; DataOut466  <=  DataIn2; DataOut467  <=  DataIn3; end
5  : begin DataOut468  <=  DataIn0; DataOut469  <=  DataIn1; DataOut470  <=  DataIn2; DataOut471  <=  DataIn3; end
6  : begin DataOut472  <=  DataIn0; DataOut473  <=  DataIn1; DataOut474  <=  DataIn2; DataOut475  <=  DataIn3; end
7  : begin DataOut476  <=  DataIn0; DataOut477  <=  DataIn1; DataOut478  <=  DataIn2; DataOut479  <=  DataIn3; end
8  : begin DataOut480  <=  DataIn0; DataOut481  <=  DataIn1; DataOut482  <=  DataIn2; DataOut483  <=  DataIn3; end
9  : begin DataOut484  <=  DataIn0; DataOut485  <=  DataIn1; DataOut486  <=  DataIn2; DataOut487  <=  DataIn3; end
10  : begin DataOut488  <=  DataIn0; DataOut489  <=  DataIn1; DataOut490  <=  DataIn2; DataOut491  <=  DataIn3; end
11  : begin DataOut492  <=  DataIn0; DataOut493  <=  DataIn1; DataOut494  <=  DataIn2; DataOut495  <=  DataIn3; end
12  : begin DataOut496  <=  DataIn0; DataOut497  <=  DataIn1; DataOut498  <=  DataIn2; DataOut499  <=  DataIn3; end
13  : begin DataOut500  <=  DataIn0; DataOut501  <=  DataIn1; DataOut502  <=  DataIn2; DataOut503  <=  DataIn3; end
14  : begin DataOut504  <=  DataIn0; DataOut505  <=  DataIn1; DataOut506  <=  DataIn2; DataOut507  <=  DataIn3; end
15  : begin DataOut508  <=  DataIn0; DataOut509  <=  DataIn1; DataOut510  <=  DataIn2; DataOut511  <=  DataIn3; end
16  : begin DataOut512  <=  DataIn0; DataOut513  <=  DataIn1; DataOut514  <=  DataIn2; DataOut515  <=  DataIn3; end
17  : begin DataOut516  <=  DataIn0; DataOut517  <=  DataIn1; DataOut518  <=  DataIn2; DataOut519  <=  DataIn3; end
18  : begin DataOut520  <=  DataIn0; DataOut521  <=  DataIn1; DataOut522  <=  DataIn2; DataOut523  <=  DataIn3; end
19  : begin DataOut524  <=  DataIn0; DataOut525  <=  DataIn1; DataOut526  <=  DataIn2; DataOut527  <=  DataIn3; end
20  : begin DataOut528  <=  DataIn0; DataOut529  <=  DataIn1; DataOut530  <=  DataIn2; DataOut531  <=  DataIn3; end
21  : begin DataOut532  <=  DataIn0; DataOut533  <=  DataIn1; DataOut534  <=  DataIn2; DataOut535  <=  DataIn3; end
22  : begin DataOut536  <=  DataIn0; DataOut537  <=  DataIn1; DataOut538  <=  DataIn2; DataOut539  <=  DataIn3; end
23  : begin DataOut540  <=  DataIn0; DataOut541  <=  DataIn1; DataOut542  <=  DataIn2; DataOut543  <=  DataIn3; end
24  : begin DataOut544  <=  DataIn0; DataOut545  <=  DataIn1; DataOut546  <=  DataIn2; DataOut547  <=  DataIn3; end
25  : begin DataOut548  <=  DataIn0; DataOut549  <=  DataIn1; DataOut550  <=  DataIn2; DataOut551  <=  DataIn3; end
26  : begin DataOut552  <=  DataIn0; DataOut553  <=  DataIn1; DataOut554  <=  DataIn2; DataOut555  <=  DataIn3; end
27  : begin DataOut556  <=  DataIn0; DataOut557  <=  DataIn1; DataOut558  <=  DataIn2; DataOut559  <=  DataIn3; end
28  : begin DataOut560  <=  DataIn0; DataOut561  <=  DataIn1; DataOut562  <=  DataIn2; DataOut563  <=  DataIn3; end
29  : begin DataOut564  <=  DataIn0; DataOut565  <=  DataIn1; DataOut566  <=  DataIn2; DataOut567  <=  DataIn3; end
30  : begin DataOut568  <=  DataIn0; DataOut569  <=  DataIn1; DataOut570  <=  DataIn2; DataOut571  <=  DataIn3; end
31  : begin DataOut572  <=  DataIn0; DataOut573  <=  DataIn1; DataOut574  <=  DataIn2; DataOut575  <=  DataIn3; end
32  : begin DataOut576  <=  DataIn0; DataOut577  <=  DataIn1; DataOut578  <=  DataIn2; DataOut579  <=  DataIn3; end
33  : begin DataOut580  <=  DataIn0; DataOut581  <=  DataIn1; DataOut582  <=  DataIn2; DataOut583  <=  DataIn3; end
34  : begin DataOut584  <=  DataIn0; DataOut585  <=  DataIn1; DataOut586  <=  DataIn2; DataOut587  <=  DataIn3; end
35  : begin DataOut588  <=  DataIn0; DataOut589  <=  DataIn1; DataOut590  <=  DataIn2; DataOut591  <=  DataIn3; end
36  : begin DataOut592  <=  DataIn0; DataOut593  <=  DataIn1; DataOut594  <=  DataIn2; DataOut595  <=  DataIn3; end
37  : begin DataOut596  <=  DataIn0; DataOut597  <=  DataIn1; DataOut598  <=  DataIn2; DataOut599  <=  DataIn3; end
38  : begin DataOut600  <=  DataIn0; DataOut601  <=  DataIn1; DataOut602  <=  DataIn2; DataOut603  <=  DataIn3; end
39  : begin DataOut604  <=  DataIn0; DataOut605  <=  DataIn1; DataOut606  <=  DataIn2; DataOut607  <=  DataIn3; end
40  : begin DataOut608  <=  DataIn0; DataOut609  <=  DataIn1; DataOut610  <=  DataIn2; DataOut611  <=  DataIn3; end
41  : begin DataOut612  <=  DataIn0; DataOut613  <=  DataIn1; DataOut614  <=  DataIn2; DataOut615  <=  DataIn3; end
42  : begin DataOut616  <=  DataIn0; DataOut617  <=  DataIn1; DataOut618  <=  DataIn2; DataOut619  <=  DataIn3; end
43  : begin DataOut620  <=  DataIn0; DataOut621  <=  DataIn1; DataOut622  <=  DataIn2; DataOut623  <=  DataIn3; end
44  : begin DataOut624  <=  DataIn0; DataOut625  <=  DataIn1; DataOut626  <=  DataIn2; DataOut627  <=  DataIn3; end
45  : begin DataOut628  <=  DataIn0; DataOut629  <=  DataIn1; DataOut630  <=  DataIn2; DataOut631  <=  DataIn3; end
46  : begin DataOut632  <=  DataIn0; DataOut633  <=  DataIn1; DataOut634  <=  DataIn2; DataOut635  <=  DataIn3; end
47  : begin DataOut636  <=  DataIn0; DataOut637  <=  DataIn1; DataOut638  <=  DataIn2; DataOut639  <=  DataIn3; end
48  : begin DataOut640  <=  DataIn0; DataOut641  <=  DataIn1; DataOut642  <=  DataIn2; DataOut643  <=  DataIn3; end
49  : begin DataOut644  <=  DataIn0; DataOut645  <=  DataIn1; DataOut646  <=  DataIn2; DataOut647  <=  DataIn3; end
50  : begin DataOut648  <=  DataIn0; DataOut649  <=  DataIn1; DataOut650  <=  DataIn2; DataOut651  <=  DataIn3; end
51  : begin DataOut652  <=  DataIn0; DataOut653  <=  DataIn1; DataOut654  <=  DataIn2; DataOut655  <=  DataIn3; end
52  : begin DataOut656  <=  DataIn0; DataOut657  <=  DataIn1; DataOut658  <=  DataIn2; DataOut659  <=  DataIn3; end
53  : begin DataOut660  <=  DataIn0; DataOut661  <=  DataIn1; DataOut662  <=  DataIn2; DataOut663  <=  DataIn3; end
54  : begin DataOut664  <=  DataIn0; DataOut665  <=  DataIn1; DataOut666  <=  DataIn2; DataOut667  <=  DataIn3; end
55  : begin DataOut668  <=  DataIn0; DataOut669  <=  DataIn1; DataOut670  <=  DataIn2; DataOut671  <=  DataIn3; end
56  : begin DataOut672  <=  DataIn0; DataOut673  <=  DataIn1; DataOut674  <=  DataIn2; DataOut675  <=  DataIn3; end
57  : begin DataOut676  <=  DataIn0; DataOut677  <=  DataIn1; DataOut678  <=  DataIn2; DataOut679  <=  DataIn3; end
58  : begin DataOut680  <=  DataIn0; DataOut681  <=  DataIn1; DataOut682  <=  DataIn2; DataOut683  <=  DataIn3; end
59  : begin DataOut684  <=  DataIn0; DataOut685  <=  DataIn1; DataOut686  <=  DataIn2; DataOut687  <=  DataIn3; end
60  : begin DataOut688  <=  DataIn0; DataOut689  <=  DataIn1; DataOut690  <=  DataIn2; DataOut691  <=  DataIn3; end
61  : begin DataOut692  <=  DataIn0; DataOut693  <=  DataIn1; DataOut694  <=  DataIn2; DataOut695  <=  DataIn3; end
62  : begin DataOut696  <=  DataIn0; DataOut697  <=  DataIn1; DataOut698  <=  DataIn2; DataOut699  <=  DataIn3; end
63  : begin DataOut700  <=  DataIn0; DataOut701  <=  DataIn1; DataOut702  <=  DataIn2; DataOut703  <=  DataIn3; end
64  : begin DataOut704  <=  DataIn0; DataOut705  <=  DataIn1; DataOut706  <=  DataIn2; DataOut707  <=  DataIn3; end
65  : begin DataOut708  <=  DataIn0; DataOut709  <=  DataIn1; DataOut710  <=  DataIn2; DataOut711  <=  DataIn3; end
66  : begin DataOut712  <=  DataIn0; DataOut713  <=  DataIn1; DataOut714  <=  DataIn2; DataOut715  <=  DataIn3; end
67  : begin DataOut716  <=  DataIn0; DataOut717  <=  DataIn1; DataOut718  <=  DataIn2; DataOut719  <=  DataIn3; end
68  : begin DataOut720  <=  DataIn0; DataOut721  <=  DataIn1; DataOut722  <=  DataIn2; DataOut723  <=  DataIn3; end
69  : begin DataOut724  <=  DataIn0; DataOut725  <=  DataIn1; DataOut726  <=  DataIn2; DataOut727  <=  DataIn3; end
70  : begin DataOut728  <=  DataIn0; DataOut729  <=  DataIn1; DataOut730  <=  DataIn2; DataOut731  <=  DataIn3; end
71  : begin DataOut732  <=  DataIn0; DataOut733  <=  DataIn1; DataOut734  <=  DataIn2; DataOut735  <=  DataIn3; end
72  : begin DataOut736  <=  DataIn0; DataOut737  <=  DataIn1; DataOut738  <=  DataIn2; DataOut739  <=  DataIn3; end
73  : begin DataOut740  <=  DataIn0; DataOut741  <=  DataIn1; DataOut742  <=  DataIn2; DataOut743  <=  DataIn3; end
74  : begin DataOut744  <=  DataIn0; DataOut745  <=  DataIn1; DataOut746  <=  DataIn2; DataOut747  <=  DataIn3; end
75  : begin DataOut748  <=  DataIn0; DataOut749  <=  DataIn1; DataOut750  <=  DataIn2; DataOut751  <=  DataIn3; end
76  : begin DataOut752  <=  DataIn0; DataOut753  <=  DataIn1; DataOut754  <=  DataIn2; DataOut755  <=  DataIn3; end
77  : begin DataOut756  <=  DataIn0; DataOut757  <=  DataIn1; DataOut758  <=  DataIn2; DataOut759  <=  DataIn3; end
78  : begin DataOut760  <=  DataIn0; DataOut761  <=  DataIn1; DataOut762  <=  DataIn2; DataOut763  <=  DataIn3; end
79  : begin DataOut764  <=  DataIn0; DataOut765  <=  DataIn1; DataOut766  <=  DataIn2; DataOut767  <=  DataIn3; end
80  : begin DataOut768  <=  DataIn0; DataOut769  <=  DataIn1; DataOut770  <=  DataIn2; DataOut771  <=  DataIn3; end
81  : begin DataOut772  <=  DataIn0; DataOut773  <=  DataIn1; DataOut774  <=  DataIn2; DataOut775  <=  DataIn3; end
82  : begin DataOut776  <=  DataIn0; DataOut777  <=  DataIn1; DataOut778  <=  DataIn2; DataOut779  <=  DataIn3; end
83  : begin DataOut780  <=  DataIn0; DataOut781  <=  DataIn1; DataOut782  <=  DataIn2; DataOut783  <=  DataIn3; end
84  : begin L0FINISH<= 1; end //$display("four");
default: begin L0FINISH<= 1; end //$display("five");


endcase
end
 //$display("six"); 
end

endmodule


