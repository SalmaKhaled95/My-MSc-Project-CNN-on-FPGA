//line 1
module CONV2_main_fsm (clk, rst, counter, address);
input clk,rst;
input [7:0] counter;
output reg  [3:0] address;
localparam [3:0]
W1 =4'b0 ,
W2 =4'b1 ,
W3 =4'b10 ,
W4 =4'b11 ,
W5 =4'b100 ,
W6 =4'b101 ,
W7 =4'b110 ,
W8 =4'b111 ,
W9 =4'b1000 ,
BIAS =4'b1001, WRITE =4'b1010;
reg [3:0] current_state, next_state;
always@ (counter, current_state)
begin 
case (current_state)
W1: 
 begin address=4'b0; //0
if (counter == 13) begin next_state = W2; end else begin next_state = W1; end end// i done0
W2: 
 begin address=4'b1; //1
if (counter == 26) begin next_state = W3; end else begin next_state = W2; end end// i done1
W3: 
 begin address=4'b10; //2
if (counter == 39) begin next_state = W4; end else begin next_state = W3; end end// i done2
W4: 
 begin address=4'b11; //3
if (counter == 52) begin next_state = W5; end else begin next_state = W4; end end// i done3
W5: 
 begin address=4'b100; //4
if (counter == 65) begin next_state = W6; end else begin next_state = W5; end end// i done4
W6: 
 begin address=4'b101; //5
if (counter == 78) begin next_state = W7; end else begin next_state = W6; end end// i done5
W7: 
 begin address=4'b110; //6
if (counter == 91) begin next_state = W8; end else begin next_state = W7; end end// i done6
W8: 
 begin address=4'b111; //7
if (counter == 104) begin next_state = W9; end else begin next_state = W8; end end// i done7
W9: 
 begin address=4'b1000; //8
next_state = W9; end
default:
begin 
address =4'b0;
next_state = W1;
end
endcase
end
always @(posedge clk, posedge rst)
begin 
if (rst)
current_state <= W1;
else
current_state <= next_state;
end
endmodule

//line65

module MUX5X1_13  ( In0 , In1 , In2 , In3 , In4 ,sel,out);
input [33:0] In0 , In1 , In2 , In3 , In4 ;
input [6:0] sel;
output [33:0] out;
assign out =

(sel>=0 && sel<13) ? In0:
(sel>=13 && sel<26) ? In1:
(sel>=26 && sel<39) ? In2:
(sel>=39 && sel<52) ? In3:
(sel>=52 && sel<65) ? In4:

34'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz; 
endmodule




module MUX9X1_conv2 (  In0, In1, In2, In3, In4, In5, In6, In7, In8,sel,out);
input [33:0] In0, In1, In2, In3, In4, In5, In6, In7, In8;
input [3:0] sel;
output [33:0] out;
assign out =
( ! sel[3] && ! sel[2] && ! sel[1] && ! sel[0] ) ? In0 :
( ! sel[3] && ! sel[2] && ! sel[1] &&   sel[0] ) ? In1 :
( ! sel[3] && ! sel[2] &&   sel[1] && ! sel[0] ) ? In2 :
( ! sel[3] && ! sel[2] &&   sel[1] &&   sel[0] ) ? In3 :
( ! sel[3] &&   sel[2] && ! sel[1] && ! sel[0] ) ? In4 :
( ! sel[3] &&   sel[2] && ! sel[1] &&   sel[0] ) ? In5 :
( ! sel[3] &&   sel[2] &&   sel[1] && ! sel[0] ) ? In6 :
( ! sel[3] &&   sel[2] &&   sel[1] &&   sel[0] ) ? In7 :
(   sel[3] && ! sel[2] && ! sel[1] && ! sel[0] ) ? In8 :
34'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz; 
endmodule

///////////////conv1 layer///////////////////////
//line 101

///march

module RELU(Original , clk , Modified);
input [33:0] Original;
input clk;
output reg [33:0] Modified;
always @ (posedge clk) begin 
if (Original[31]) begin Modified <=34'b0000000000000000000000000000000000; end
else begin Modified <= Original ;end
end
endmodule

//ram output
//line116
module OneRegister (clk, write, DataIn, DataOut); //ok
input clk, write;
input [33:0] DataIn;
output reg [33:0] DataOut;
initial begin DataOut <=34'b0000000000000000000000000000000000; end
always @ (posedge clk) begin 
if (write) begin DataOut <=  DataIn;  end
end
endmodule



////////////////////////////////////////////maxpool1 start //////
//line131
module COMPARATOR_MAX_TRY_tssssst( clk, A,B, C, D, Data);
input clk;

input wire [33:0] A;
input wire [33:0] B;
input wire [33:0] C;
input wire [33:0] D;

output reg [33:0] Data;

reg [33:0] AB;
reg [33:0] CD;


//initial begin $monitor("A = %b, B = %b, C = %b,  D = %b , AB = %b, CD = %b, Data= %b ",  A, B, C,  D, AB, CD, Data); end


FPComparator_8_23_F400_uid2 CompInstanceAB (clk , A , B ,  unorderedAB,  AltB , AeqB , AgtB , AleB , AgeB );
FPComparator_8_23_F400_uid2 CompInstanceCD (clk , C , D ,  unorderedCD,  CltD , CeqD , CgtD , CleD , CgeD );

always @ (posedge clk) begin
if (AltB && CltD) begin  AB = B; CD = D;  end
else if (AgeB && CltD) begin AB = A ; CD  =D  ;  end
else if (AltB && CgeD) begin  AB =  B ; CD  = C ; end
else if (AgeB && CgeD) begin AB = A ; CD  = C ;  end
end

FPComparator_8_23_F400_uid2 CompInstanceABCD (clk ,AB , CD ,  unorderedABCD,  ABltCD , ABeqCD , ABgtCD , ABleCD , ABgeCD );
always @ (posedge clk) begin
if (ABgeCD) begin  Data = AB;  end
else if (ABltCD) begin  Data = CD;  end
else begin Data = 34'b0; end
end


endmodule

//////////////////layer2 conv
///march
//line170

module OneRegister_In4_xBIAS (clk, write, DataIn, DataOut);
input clk, write; input [33:0] DataIn; output reg [33:0] DataOut;
//initial begin DataOut <= 66'b011011111110000011010101101110001100000000000000000000000000000000
initial begin DataOut <=   34'b0110111100000110101011011100011000
 ; end
always @ (posedge clk) begin if (write) begin DataOut <=  DataIn;  end end endmodule
//////


//line 183

///march

 
 module In1_ROM_9x66bit_3(clk, addr, dout); input clk; input [7:0] addr; output reg [33:0] dout;
// module In4_ROM_9x66bit_0(clk, addr, dout); input clk; input [7:0] addr; output reg [65:0] dout;
always @(posedge clk) begin case(addr)
0: dout <= 34'b0100111101001001010110100111110100
 ;13: dout <= 34'b0110111110001100010010000001101010
 ;26: dout <= 34'b0110111110101011101100010001010111
 ;39: dout <= 34'b0100111101000110101110010001110110
 ;52: dout <= 34'b0100111101101010110001010100110010
 ;65: dout <= 34'b0100111101101110001110110001100111
 ;78: dout <= 34'b0110111100100100110100010110101000
 ;91: dout <= 34'b0110111100111001000100100101111101
 ;104: dout <= 34'b0100111101111100100100101011101010
 
 ;endcase end endmodule


module In2_ROM_9x66bit_3(clk, addr, dout); input clk; input [7:0] addr; output reg [33:0] dout;
//module In4_ROM_9x66bit_1(clk, addr, dout); input clk; input [7:0] addr; output reg [65:0] dout;
always @(posedge clk) begin case(addr)

0: dout <= 34'b0100111110101011000110100001111110
 ;13: dout <= 34'b0100111100100010001000001110000010
 ;26: dout <= 34'b0110111101011110001110000001111001
 ;39: dout <= 34'b0100111110111110111001110011100110
 ;52: dout <= 34'b0100111110000111111111000111001010
 ;65: dout <= 34'b0100111100010101101001110001010101
 ;78: dout <= 34'b0100111110100000110000011111111111
 ;91: dout <= 34'b0100111101101100000011101100011011
 ;104: dout <= 34'b0110111101010000001001011010100000
 
 ;endcase end endmodule


module In3_ROM_9x66bit_3(clk, addr, dout); input clk; input [7:0] addr; output reg [33:0] dout;
//module In4_ROM_9x66bit_2(clk, addr, dout); input clk; input [7:0] addr; output reg [65:0] dout;
always @(posedge clk) begin case(addr)

0: dout <= 34'b0100111110011111001000000110011110
 ;13: dout <= 34'b0100111101110110101000100011100010
 ;26: dout <= 34'b0100111111000000011100010100010011
 ;39: dout <= 34'b0100111110101011010100101010001001
 ;52: dout <= 34'b0100111110010101000100110001110111
 ;65: dout <= 34'b0100111110010010011111001010001111
 ;78: dout <= 34'b0110111110101000010010001100100110
 ;91: dout <= 34'b0110111110001101111001100010111011
 ;104: dout <= 34'b0110111110001000011101000011000001
 
 ;endcase end endmodule

module In4_ROM_9x66bit_3(clk, addr, dout); input clk; input [7:0] addr; output reg [33:0] dout;
//module In4_ROM_9x66bit_3(clk, addr, dout); input clk; input [7:0] addr; output reg [65:0] dout;
always @(posedge clk) begin case(addr)

0: dout <= 34'b0100111110001000101010101001101101
 ;13: dout <= 34'b0110111100000111110101110011101011
 ;26: dout <= 34'b0100111111000111110101001111011110
 ;39: dout <= 34'b0110111100100011000000011000101000
 ;52: dout <= 34'b0100111101111101101101001000101001
 ;65: dout <= 34'b0100111110100110001011111001011001
 ;78: dout <= 34'b0110111110011011101000000000101000
 ;91: dout <= 34'b0110111101101110001000011111111011
 ;104: dout <= 34'b0100111100111000100011111100100010
 
 ;endcase end endmodule
 ///////
//channel 1 of all filters



//dense2
//line 247



module AXIinputFromARM_3_1(clk, AXIinput, AXIstart , L0FINISH, 
REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143 
);


input clk, AXIstart;
input [31:0] AXIinput;
output reg [33:0] REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143;
output reg [33:0] REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 ;
output reg [33:0] REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 ;
output reg [33:0] REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143;
output reg L0FINISH;


wire [10:0] counter; 
COUNTER_LAYER_1200_cycles TheCounter (clk, counter, AXIstart);
initial begin L0FINISH <= 1'b0; end
always @(posedge clk) 
begin 
if (AXIstart && !L0FINISH)
begin

case(counter) 

0  : begin {REGofMAX1DataOut_F1_0[33:2] } <= AXIinput ; end 
1  : begin {REGofMAX1DataOut_F1_0[1:0] , REGofMAX1DataOut_F1_1[33:4] } <= AXIinput ; end 
2  : begin {REGofMAX1DataOut_F1_1[3:0] , REGofMAX1DataOut_F1_2[33:6]  } <= AXIinput ; end 
3  : begin {REGofMAX1DataOut_F1_2[5:0] , REGofMAX1DataOut_F1_3[33:8]  } <= AXIinput ; end 
4  : begin {REGofMAX1DataOut_F1_3[7:0] , REGofMAX1DataOut_F1_4[33:10]  } <= AXIinput ; end 
5  : begin {REGofMAX1DataOut_F1_4[9:0] , REGofMAX1DataOut_F1_5[33:12]  } <= AXIinput ; end 
6  : begin {REGofMAX1DataOut_F1_5[11:0] , REGofMAX1DataOut_F1_6[33:14] } <= AXIinput ; end 
7  : begin {REGofMAX1DataOut_F1_6[13:0] , REGofMAX1DataOut_F1_7[33:16] } <= AXIinput ; end 
8  : begin {REGofMAX1DataOut_F1_7[15:0] , REGofMAX1DataOut_F1_8[33:18] } <= AXIinput ; end 
9  : begin {REGofMAX1DataOut_F1_8[17:0] , REGofMAX1DataOut_F1_9[33:20] } <= AXIinput ; end 
10  : begin {REGofMAX1DataOut_F1_9[19:0] , REGofMAX1DataOut_F1_10[33:22] } <= AXIinput ; end 
11  : begin {REGofMAX1DataOut_F1_10[21:0] , REGofMAX1DataOut_F1_11[33:24] } <= AXIinput ; end  
12  : begin {REGofMAX1DataOut_F1_11[23:0] , REGofMAX1DataOut_F1_12[33:26] } <= AXIinput ; end 
13  : begin {REGofMAX1DataOut_F1_12[25:0] , REGofMAX1DataOut_F1_13[33:28] } <= AXIinput ; end 
14  : begin {REGofMAX1DataOut_F1_13[27:0] , REGofMAX1DataOut_F1_14[33:30] } <= AXIinput ; end 
15  : begin {REGofMAX1DataOut_F1_14[29:0] , REGofMAX1DataOut_F1_15[33:32] } <= AXIinput ; end 
16  : begin {REGofMAX1DataOut_F1_15[31:0] } <= AXIinput ; end 
17  : begin {REGofMAX1DataOut_F1_16[33:2] } <= AXIinput ; end 
18  : begin {REGofMAX1DataOut_F1_16[1:0], REGofMAX1DataOut_F1_17[33:4] } <= AXIinput ; end 
19  : begin {REGofMAX1DataOut_F1_17[3:0] , REGofMAX1DataOut_F1_18[33:6]  } <= AXIinput ; end 
20  : begin {REGofMAX1DataOut_F1_18[5:0] , REGofMAX1DataOut_F1_19[33:8]  } <= AXIinput ; end 
21  : begin {REGofMAX1DataOut_F1_19[7:0] , REGofMAX1DataOut_F1_20[33:10]  } <= AXIinput ; end 
22  : begin {REGofMAX1DataOut_F1_20[9:0] , REGofMAX1DataOut_F1_21[33:12]  } <= AXIinput ; end 
23  : begin {REGofMAX1DataOut_F1_21[11:0] , REGofMAX1DataOut_F1_22[33:14] } <= AXIinput ; end 
24  : begin {REGofMAX1DataOut_F1_22[13:0] , REGofMAX1DataOut_F1_23[33:16] } <= AXIinput ; end 
25  : begin {REGofMAX1DataOut_F1_23[15:0] , REGofMAX1DataOut_F1_24[33:18] } <= AXIinput ; end 
26  : begin {REGofMAX1DataOut_F1_24[17:0] , REGofMAX1DataOut_F1_25[33:20] } <= AXIinput ; end 
27  : begin {REGofMAX1DataOut_F1_25[19:0] , REGofMAX1DataOut_F1_26[33:22] } <= AXIinput ; end 
28  : begin {REGofMAX1DataOut_F1_26[21:0] , REGofMAX1DataOut_F1_27[33:24] } <= AXIinput ; end  
29  : begin {REGofMAX1DataOut_F1_27[23:0] , REGofMAX1DataOut_F1_28[33:26] } <= AXIinput ; end 
30  : begin {REGofMAX1DataOut_F1_28[25:0] , REGofMAX1DataOut_F1_29[33:28] } <= AXIinput ; end 
31  : begin {REGofMAX1DataOut_F1_29[27:0] , REGofMAX1DataOut_F1_30[33:30] } <= AXIinput ; end 
32  : begin {REGofMAX1DataOut_F1_30[29:0] , REGofMAX1DataOut_F1_31[33:32] } <= AXIinput ; end 
33  : begin {REGofMAX1DataOut_F1_31[31:0] } <= AXIinput ; end 
34  : begin {REGofMAX1DataOut_F1_32[33:2] } <= AXIinput ; end 
35  : begin {REGofMAX1DataOut_F1_32[1:0], REGofMAX1DataOut_F1_33[33:4] } <= AXIinput ; end 
36  : begin {REGofMAX1DataOut_F1_33[3:0] , REGofMAX1DataOut_F1_34[33:6]  } <= AXIinput ; end 
37  : begin {REGofMAX1DataOut_F1_34[5:0] , REGofMAX1DataOut_F1_35[33:8]  } <= AXIinput ; end 
38  : begin {REGofMAX1DataOut_F1_35[7:0] , REGofMAX1DataOut_F1_36[33:10]  } <= AXIinput ; end 
39  : begin {REGofMAX1DataOut_F1_36[9:0] , REGofMAX1DataOut_F1_37[33:12]  } <= AXIinput ; end 
40  : begin {REGofMAX1DataOut_F1_37[11:0] , REGofMAX1DataOut_F1_38[33:14] } <= AXIinput ; end  
41  : begin {REGofMAX1DataOut_F1_38[13:0] , REGofMAX1DataOut_F1_39[33:16] } <= AXIinput ; end 
42  : begin {REGofMAX1DataOut_F1_39[15:0] , REGofMAX1DataOut_F1_40[33:18] } <= AXIinput ; end 
43  : begin {REGofMAX1DataOut_F1_40[17:0] , REGofMAX1DataOut_F1_41[33:20] } <= AXIinput ; end 
44  : begin {REGofMAX1DataOut_F1_41[19:0] , REGofMAX1DataOut_F1_42[33:22] } <= AXIinput ; end  
45  : begin {REGofMAX1DataOut_F1_42[21:0] , REGofMAX1DataOut_F1_43[33:24] } <= AXIinput ; end 
46  : begin {REGofMAX1DataOut_F1_43[23:0] , REGofMAX1DataOut_F1_44[33:26] } <= AXIinput ; end 
47  : begin {REGofMAX1DataOut_F1_44[25:0] , REGofMAX1DataOut_F1_45[33:28] } <= AXIinput ; end  
48  : begin {REGofMAX1DataOut_F1_45[27:0] , REGofMAX1DataOut_F1_46[33:30] } <= AXIinput ; end 
49  : begin {REGofMAX1DataOut_F1_46[29:0] , REGofMAX1DataOut_F1_47[33:32] } <= AXIinput ; end 
50  : begin {REGofMAX1DataOut_F1_47[31:0] } <= AXIinput ; end
51  : begin {REGofMAX1DataOut_F1_48[33:2] } <= AXIinput ; end 
52  : begin {REGofMAX1DataOut_F1_48[1:0], REGofMAX1DataOut_F1_49[33:4] } <= AXIinput ; end 
53  : begin {REGofMAX1DataOut_F1_49[3:0] , REGofMAX1DataOut_F1_50[33:6]  } <= AXIinput ; end 
54  : begin {REGofMAX1DataOut_F1_50[5:0] , REGofMAX1DataOut_F1_51[33:8]  } <= AXIinput ; end 
55  : begin {REGofMAX1DataOut_F1_51[7:0] , REGofMAX1DataOut_F1_52[33:10]  } <= AXIinput ; end 
56  : begin {REGofMAX1DataOut_F1_52[9:0] , REGofMAX1DataOut_F1_53[33:12]  } <= AXIinput ; end 
57  : begin {REGofMAX1DataOut_F1_53[11:0] , REGofMAX1DataOut_F1_54[33:14] } <= AXIinput ; end 
58  : begin {REGofMAX1DataOut_F1_54[13:0] , REGofMAX1DataOut_F1_55[33:16] } <= AXIinput ; end 
59  : begin {REGofMAX1DataOut_F1_55[15:0] , REGofMAX1DataOut_F1_56[33:18] } <= AXIinput ; end 
60  : begin {REGofMAX1DataOut_F1_56[17:0] , REGofMAX1DataOut_F1_57[33:20] } <= AXIinput ; end 
61  : begin {REGofMAX1DataOut_F1_57[19:0] , REGofMAX1DataOut_F1_58[33:22] } <= AXIinput ; end 
62  : begin {REGofMAX1DataOut_F1_58[21:0] , REGofMAX1DataOut_F1_59[33:24] } <= AXIinput ; end 
63  : begin {REGofMAX1DataOut_F1_59[23:0] , REGofMAX1DataOut_F1_60[33:26] } <= AXIinput ; end  
64  : begin {REGofMAX1DataOut_F1_60[25:0] , REGofMAX1DataOut_F1_61[33:28] } <= AXIinput ; end  
65  : begin {REGofMAX1DataOut_F1_61[27:0] , REGofMAX1DataOut_F1_62[33:30] } <= AXIinput ; end 
66 : begin {REGofMAX1DataOut_F1_62[29:0] , REGofMAX1DataOut_F1_63[33:32] } <= AXIinput ; end 
67  : begin {REGofMAX1DataOut_F1_63[31:0] } <= AXIinput ; end 
68  : begin {REGofMAX1DataOut_F1_64[33:2] } <= AXIinput ; end 
69  : begin {REGofMAX1DataOut_F1_64[1:0], REGofMAX1DataOut_F1_65[33:4] } <= AXIinput ; end 
70  : begin {REGofMAX1DataOut_F1_65[3:0] , REGofMAX1DataOut_F1_66[33:6]  } <= AXIinput ; end  
71  : begin {REGofMAX1DataOut_F1_66[5:0] , REGofMAX1DataOut_F1_67[33:8]  } <= AXIinput ; end 
72  : begin {REGofMAX1DataOut_F1_67[7:0] , REGofMAX1DataOut_F1_68[33:10]  } <= AXIinput ; end 
73  : begin {REGofMAX1DataOut_F1_68[9:0] , REGofMAX1DataOut_F1_69[33:12]  } <= AXIinput ; end 
74  : begin {REGofMAX1DataOut_F1_69[11:0] , REGofMAX1DataOut_F1_70[33:14] } <= AXIinput ; end 
75  : begin {REGofMAX1DataOut_F1_70[13:0] , REGofMAX1DataOut_F1_71[33:16] } <= AXIinput ; end 
76  : begin {REGofMAX1DataOut_F1_71[15:0] , REGofMAX1DataOut_F1_72[33:18] } <= AXIinput ; end  
77  : begin {REGofMAX1DataOut_F1_72[17:0] , REGofMAX1DataOut_F1_73[33:20] } <= AXIinput ; end 
78  : begin {REGofMAX1DataOut_F1_73[19:0] , REGofMAX1DataOut_F1_74[33:22] } <= AXIinput ; end 
79  : begin {REGofMAX1DataOut_F1_74[21:0] , REGofMAX1DataOut_F1_75[33:24] } <= AXIinput ; end 
80  : begin {REGofMAX1DataOut_F1_75[23:0] , REGofMAX1DataOut_F1_76[33:26] } <= AXIinput ; end 
81  : begin {REGofMAX1DataOut_F1_76[25:0] , REGofMAX1DataOut_F1_77[33:28] } <= AXIinput ; end 
82  : begin {REGofMAX1DataOut_F1_77[27:0] , REGofMAX1DataOut_F1_78[33:30] } <= AXIinput ; end 
83  : begin {REGofMAX1DataOut_F1_78[29:0] , REGofMAX1DataOut_F1_79[33:32] } <= AXIinput ; end 
84  : begin {REGofMAX1DataOut_F1_79[31:0] } <= AXIinput ; end 
85  : begin {REGofMAX1DataOut_F1_80[33:2] } <= AXIinput ; end 
86  : begin {REGofMAX1DataOut_F1_80[1:0], REGofMAX1DataOut_F1_81[33:4] } <= AXIinput ; end 
87  : begin {REGofMAX1DataOut_F1_81[3:0] , REGofMAX1DataOut_F1_82[33:6]  } <= AXIinput ; end 
88  : begin {REGofMAX1DataOut_F1_82[5:0] , REGofMAX1DataOut_F1_83[33:8]  } <= AXIinput ; end 
89  : begin {REGofMAX1DataOut_F1_83[7:0] , REGofMAX1DataOut_F1_84[33:10]  } <= AXIinput ; end 
90  : begin {REGofMAX1DataOut_F1_84[9:0] , REGofMAX1DataOut_F1_85[33:12]  } <= AXIinput ; end 
91  : begin {REGofMAX1DataOut_F1_85[11:0] , REGofMAX1DataOut_F1_86[33:14] } <= AXIinput ; end  
92  : begin {REGofMAX1DataOut_F1_86[13:0] , REGofMAX1DataOut_F1_87[33:16] } <= AXIinput ; end 
93  : begin {REGofMAX1DataOut_F1_87[15:0] , REGofMAX1DataOut_F1_88[33:18] } <= AXIinput ; end 
94  : begin {REGofMAX1DataOut_F1_88[17:0] , REGofMAX1DataOut_F1_89[33:20] } <= AXIinput ; end 
95  : begin {REGofMAX1DataOut_F1_89[19:0] , REGofMAX1DataOut_F1_90[33:22] } <= AXIinput ; end 
96  : begin {REGofMAX1DataOut_F1_90[21:0] , REGofMAX1DataOut_F1_91[33:24] } <= AXIinput ; end 
97  : begin {REGofMAX1DataOut_F1_91[23:0] , REGofMAX1DataOut_F1_92[33:26] } <= AXIinput ; end 
98  : begin {REGofMAX1DataOut_F1_92[25:0] , REGofMAX1DataOut_F1_93[33:28] } <= AXIinput ; end 
99  : begin {REGofMAX1DataOut_F1_93[27:0] , REGofMAX1DataOut_F1_94[33:30] } <= AXIinput ; end 
100  : begin {REGofMAX1DataOut_F1_94[29:0] , REGofMAX1DataOut_F1_95[33:32] } <= AXIinput ; end 
101  : begin {REGofMAX1DataOut_F1_95[31:0] } <= AXIinput ; end 
102  : begin {REGofMAX1DataOut_F1_96[33:2] } <= AXIinput ; end 
103  : begin {REGofMAX1DataOut_F1_96[1:0], REGofMAX1DataOut_F1_97[33:4] } <= AXIinput ; end 
104  : begin {REGofMAX1DataOut_F1_97[3:0] , REGofMAX1DataOut_F1_98[33:6]  } <= AXIinput ; end 
105  : begin {REGofMAX1DataOut_F1_98[5:0] , REGofMAX1DataOut_F1_99[33:8]  } <= AXIinput ; end  
106  : begin {REGofMAX1DataOut_F1_99[7:0] , REGofMAX1DataOut_F1_100[33:10]  } <= AXIinput ; end 
107  : begin {REGofMAX1DataOut_F1_100[9:0] , REGofMAX1DataOut_F1_101[33:12]  } <= AXIinput ; end 
108  : begin {REGofMAX1DataOut_F1_101[11:0] , REGofMAX1DataOut_F1_102[33:14] } <= AXIinput ; end  
109  : begin {REGofMAX1DataOut_F1_102[13:0] , REGofMAX1DataOut_F1_103[33:16] } <= AXIinput ; end 
110  : begin {REGofMAX1DataOut_F1_103[15:0] , REGofMAX1DataOut_F1_104[33:18] } <= AXIinput ; end 
111  : begin {REGofMAX1DataOut_F1_104[17:0] , REGofMAX1DataOut_F1_105[33:20] } <= AXIinput ; end 
112  : begin {REGofMAX1DataOut_F1_105[19:0] , REGofMAX1DataOut_F1_106[33:22] } <= AXIinput ; end 
113  : begin {REGofMAX1DataOut_F1_106[21:0] , REGofMAX1DataOut_F1_107[33:24] } <= AXIinput ; end 
114  : begin {REGofMAX1DataOut_F1_107[23:0] , REGofMAX1DataOut_F1_108[33:26] } <= AXIinput ; end 
115  : begin {REGofMAX1DataOut_F1_108[25:0] , REGofMAX1DataOut_F1_109[33:28] } <= AXIinput ; end 
116  : begin {REGofMAX1DataOut_F1_109[27:0] , REGofMAX1DataOut_F1_110[33:30] } <= AXIinput ; end 
117  : begin {REGofMAX1DataOut_F1_110[29:0] , REGofMAX1DataOut_F1_111[33:32] } <= AXIinput ; end 
118  : begin {REGofMAX1DataOut_F1_111[31:0] } <= AXIinput ; end 
119  : begin {REGofMAX1DataOut_F1_112[33:2] } <= AXIinput ; end 
120  : begin {REGofMAX1DataOut_F1_112[1:0], REGofMAX1DataOut_F1_113[33:4] } <= AXIinput ; end 
121  : begin {REGofMAX1DataOut_F1_113[3:0] , REGofMAX1DataOut_F1_114[33:6]  } <= AXIinput ; end 
122  : begin {REGofMAX1DataOut_F1_114[5:0] , REGofMAX1DataOut_F1_115[33:8]  } <= AXIinput ; end 
123  : begin {REGofMAX1DataOut_F1_115[7:0] , REGofMAX1DataOut_F1_116[33:10]  } <= AXIinput ; end 
124  : begin {REGofMAX1DataOut_F1_116[9:0] , REGofMAX1DataOut_F1_117[33:12]  } <= AXIinput ; end 
125  : begin {REGofMAX1DataOut_F1_117[11:0] , REGofMAX1DataOut_F1_118[33:14] } <= AXIinput ; end 
126  : begin {REGofMAX1DataOut_F1_118[13:0] , REGofMAX1DataOut_F1_119[33:16] } <= AXIinput ; end 
127  : begin {REGofMAX1DataOut_F1_119[15:0] , REGofMAX1DataOut_F1_120[33:18] } <= AXIinput ; end 
128  : begin {REGofMAX1DataOut_F1_120[17:0] , REGofMAX1DataOut_F1_121[33:20] } <= AXIinput ; end 
129  : begin {REGofMAX1DataOut_F1_121[19:0] , REGofMAX1DataOut_F1_122[33:22] } <= AXIinput ; end 
130  : begin {REGofMAX1DataOut_F1_122[21:0] , REGofMAX1DataOut_F1_123[33:24] } <= AXIinput ; end 
131  : begin {REGofMAX1DataOut_F1_123[23:0] , REGofMAX1DataOut_F1_124[33:26] } <= AXIinput ; end 
132  : begin {REGofMAX1DataOut_F1_124[25:0] , REGofMAX1DataOut_F1_125[33:28] } <= AXIinput ; end 
133  : begin {REGofMAX1DataOut_F1_125[27:0] , REGofMAX1DataOut_F1_126[33:30] } <= AXIinput ; end 
134  : begin {REGofMAX1DataOut_F1_126[29:0] , REGofMAX1DataOut_F1_127[33:32] } <= AXIinput ; end 
135  : begin {REGofMAX1DataOut_F1_127[31:0] } <= AXIinput ; end 
136  : begin {REGofMAX1DataOut_F1_128[33:2] } <= AXIinput ; end 
137  : begin {REGofMAX1DataOut_F1_128[1:0], REGofMAX1DataOut_F1_129[33:4] } <= AXIinput ; end 
138  : begin {REGofMAX1DataOut_F1_129[3:0] , REGofMAX1DataOut_F1_130[33:6]  } <= AXIinput ; end 
139  : begin {REGofMAX1DataOut_F1_130[5:0] , REGofMAX1DataOut_F1_131[33:8]  } <= AXIinput ; end 
140  : begin {REGofMAX1DataOut_F1_131[7:0] , REGofMAX1DataOut_F1_132[33:10]  } <= AXIinput ; end 
141  : begin {REGofMAX1DataOut_F1_132[9:0] , REGofMAX1DataOut_F1_133[33:12]  } <= AXIinput ; end 
142  : begin {REGofMAX1DataOut_F1_133[11:0] , REGofMAX1DataOut_F1_134[33:14] } <= AXIinput ; end 
143  : begin {REGofMAX1DataOut_F1_134[13:0] , REGofMAX1DataOut_F1_135[33:16] } <= AXIinput ; end 
144  : begin {REGofMAX1DataOut_F1_135[15:0] , REGofMAX1DataOut_F1_136[33:18] } <= AXIinput ; end 
145  : begin {REGofMAX1DataOut_F1_136[17:0] , REGofMAX1DataOut_F1_137[33:20] } <= AXIinput ; end 
146  : begin {REGofMAX1DataOut_F1_137[19:0] , REGofMAX1DataOut_F1_138[33:22] } <= AXIinput ; end 
147  : begin {REGofMAX1DataOut_F1_138[21:0] , REGofMAX1DataOut_F1_139[33:24] } <= AXIinput ; end 
148  : begin {REGofMAX1DataOut_F1_139[23:0] , REGofMAX1DataOut_F1_140[33:26] } <= AXIinput ; end 
149  : begin {REGofMAX1DataOut_F1_140[25:0] , REGofMAX1DataOut_F1_141[33:28] } <= AXIinput ; end 
150  : begin {REGofMAX1DataOut_F1_141[27:0] , REGofMAX1DataOut_F1_142[33:30] } <= AXIinput ; end 
151  : begin {REGofMAX1DataOut_F1_142[29:0] , REGofMAX1DataOut_F1_143[33:32] } <= AXIinput ; end 
152  : begin {REGofMAX1DataOut_F1_143[31:0] } <= AXIinput ; end 

0  + 153 : begin {REGofMAX1DataOut_F2_0[33:2] } <= AXIinput ; end 
1  + 153 : begin {REGofMAX1DataOut_F2_0[1:0] , REGofMAX1DataOut_F2_1[33:4] } <= AXIinput ; end 
2  + 153 : begin {REGofMAX1DataOut_F2_1[3:0] , REGofMAX1DataOut_F2_2[33:6]  } <= AXIinput ; end 
3  + 153 : begin {REGofMAX1DataOut_F2_2[5:0] , REGofMAX1DataOut_F2_3[33:8]  } <= AXIinput ; end 
4  + 153 : begin {REGofMAX1DataOut_F2_3[7:0] , REGofMAX1DataOut_F2_4[33:10]  } <= AXIinput ; end 
5  + 153 : begin {REGofMAX1DataOut_F2_4[9:0] , REGofMAX1DataOut_F2_5[33:12]  } <= AXIinput ; end 
6  + 153 : begin {REGofMAX1DataOut_F2_5[11:0] , REGofMAX1DataOut_F2_6[33:14] } <= AXIinput ; end 
7  + 153 : begin {REGofMAX1DataOut_F2_6[13:0] , REGofMAX1DataOut_F2_7[33:16] } <= AXIinput ; end 
8  + 153 : begin {REGofMAX1DataOut_F2_7[15:0] , REGofMAX1DataOut_F2_8[33:18] } <= AXIinput ; end 
9  + 153 : begin {REGofMAX1DataOut_F2_8[17:0] , REGofMAX1DataOut_F2_9[33:20] } <= AXIinput ; end 
10  + 153 : begin {REGofMAX1DataOut_F2_9[19:0] , REGofMAX1DataOut_F2_10[33:22] } <= AXIinput ; end 
11  + 153 : begin {REGofMAX1DataOut_F2_10[21:0] , REGofMAX1DataOut_F2_11[33:24] } <= AXIinput ; end  
12  + 153 : begin {REGofMAX1DataOut_F2_11[23:0] , REGofMAX1DataOut_F2_12[33:26] } <= AXIinput ; end 
13  + 153 : begin {REGofMAX1DataOut_F2_12[25:0] , REGofMAX1DataOut_F2_13[33:28] } <= AXIinput ; end 
14  + 153 : begin {REGofMAX1DataOut_F2_13[27:0] , REGofMAX1DataOut_F2_14[33:30] } <= AXIinput ; end 
15  + 153 : begin {REGofMAX1DataOut_F2_14[29:0] , REGofMAX1DataOut_F2_15[33:32] } <= AXIinput ; end 
16  + 153 : begin {REGofMAX1DataOut_F2_15[31:0] } <= AXIinput ; end 
17  + 153 : begin {REGofMAX1DataOut_F2_16[33:2] } <= AXIinput ; end 
18  + 153 : begin {REGofMAX1DataOut_F2_16[1:0], REGofMAX1DataOut_F2_17[33:4] } <= AXIinput ; end 
19  + 153 : begin {REGofMAX1DataOut_F2_17[3:0] , REGofMAX1DataOut_F2_18[33:6]  } <= AXIinput ; end 
20  + 153 : begin {REGofMAX1DataOut_F2_18[5:0] , REGofMAX1DataOut_F2_19[33:8]  } <= AXIinput ; end 
21  + 153 : begin {REGofMAX1DataOut_F2_19[7:0] , REGofMAX1DataOut_F2_20[33:10]  } <= AXIinput ; end 
22  + 153 : begin {REGofMAX1DataOut_F2_20[9:0] , REGofMAX1DataOut_F2_21[33:12]  } <= AXIinput ; end 
23  + 153 : begin {REGofMAX1DataOut_F2_21[11:0] , REGofMAX1DataOut_F2_22[33:14] } <= AXIinput ; end 
24  + 153 : begin {REGofMAX1DataOut_F2_22[13:0] , REGofMAX1DataOut_F2_23[33:16] } <= AXIinput ; end 
25  + 153 : begin {REGofMAX1DataOut_F2_23[15:0] , REGofMAX1DataOut_F2_24[33:18] } <= AXIinput ; end 
26  + 153 : begin {REGofMAX1DataOut_F2_24[17:0] , REGofMAX1DataOut_F2_25[33:20] } <= AXIinput ; end 
27  + 153 : begin {REGofMAX1DataOut_F2_25[19:0] , REGofMAX1DataOut_F2_26[33:22] } <= AXIinput ; end 
28  + 153 : begin {REGofMAX1DataOut_F2_26[21:0] , REGofMAX1DataOut_F2_27[33:24] } <= AXIinput ; end  
29  + 153 : begin {REGofMAX1DataOut_F2_27[23:0] , REGofMAX1DataOut_F2_28[33:26] } <= AXIinput ; end 
30  + 153 : begin {REGofMAX1DataOut_F2_28[25:0] , REGofMAX1DataOut_F2_29[33:28] } <= AXIinput ; end 
31  + 153 : begin {REGofMAX1DataOut_F2_29[27:0] , REGofMAX1DataOut_F2_30[33:30] } <= AXIinput ; end 
32  + 153 : begin {REGofMAX1DataOut_F2_30[29:0] , REGofMAX1DataOut_F2_31[33:32] } <= AXIinput ; end 
33  + 153 : begin {REGofMAX1DataOut_F2_31[31:0] } <= AXIinput ; end 
34  + 153 : begin {REGofMAX1DataOut_F2_32[33:2] } <= AXIinput ; end 
35  + 153 : begin {REGofMAX1DataOut_F2_32[1:0], REGofMAX1DataOut_F2_33[33:4] } <= AXIinput ; end 
36  + 153 : begin {REGofMAX1DataOut_F2_33[3:0] , REGofMAX1DataOut_F2_34[33:6]  } <= AXIinput ; end 
37  + 153 : begin {REGofMAX1DataOut_F2_34[5:0] , REGofMAX1DataOut_F2_35[33:8]  } <= AXIinput ; end 
38  + 153 : begin {REGofMAX1DataOut_F2_35[7:0] , REGofMAX1DataOut_F2_36[33:10]  } <= AXIinput ; end 
39  + 153 : begin {REGofMAX1DataOut_F2_36[9:0] , REGofMAX1DataOut_F2_37[33:12]  } <= AXIinput ; end 
40  + 153 : begin {REGofMAX1DataOut_F2_37[11:0] , REGofMAX1DataOut_F2_38[33:14] } <= AXIinput ; end  
41  + 153 : begin {REGofMAX1DataOut_F2_38[13:0] , REGofMAX1DataOut_F2_39[33:16] } <= AXIinput ; end 
42  + 153 : begin {REGofMAX1DataOut_F2_39[15:0] , REGofMAX1DataOut_F2_40[33:18] } <= AXIinput ; end 
43  + 153 : begin {REGofMAX1DataOut_F2_40[17:0] , REGofMAX1DataOut_F2_41[33:20] } <= AXIinput ; end 
44  + 153 : begin {REGofMAX1DataOut_F2_41[19:0] , REGofMAX1DataOut_F2_42[33:22] } <= AXIinput ; end  
45  + 153 : begin {REGofMAX1DataOut_F2_42[21:0] , REGofMAX1DataOut_F2_43[33:24] } <= AXIinput ; end 
46  + 153 : begin {REGofMAX1DataOut_F2_43[23:0] , REGofMAX1DataOut_F2_44[33:26] } <= AXIinput ; end 
47  + 153 : begin {REGofMAX1DataOut_F2_44[25:0] , REGofMAX1DataOut_F2_45[33:28] } <= AXIinput ; end  
48  + 153 : begin {REGofMAX1DataOut_F2_45[27:0] , REGofMAX1DataOut_F2_46[33:30] } <= AXIinput ; end 
49  + 153 : begin {REGofMAX1DataOut_F2_46[29:0] , REGofMAX1DataOut_F2_47[33:32] } <= AXIinput ; end 
50  + 153 : begin {REGofMAX1DataOut_F2_47[31:0] } <= AXIinput ; end
51  + 153 : begin {REGofMAX1DataOut_F2_48[33:2] } <= AXIinput ; end 
52  + 153 : begin {REGofMAX1DataOut_F2_48[1:0], REGofMAX1DataOut_F2_49[33:4] } <= AXIinput ; end 
53  + 153 : begin {REGofMAX1DataOut_F2_49[3:0] , REGofMAX1DataOut_F2_50[33:6]  } <= AXIinput ; end 
54  + 153 : begin {REGofMAX1DataOut_F2_50[5:0] , REGofMAX1DataOut_F2_51[33:8]  } <= AXIinput ; end 
55  + 153 : begin {REGofMAX1DataOut_F2_51[7:0] , REGofMAX1DataOut_F2_52[33:10]  } <= AXIinput ; end 
56  + 153 : begin {REGofMAX1DataOut_F2_52[9:0] , REGofMAX1DataOut_F2_53[33:12]  } <= AXIinput ; end 
57  + 153 : begin {REGofMAX1DataOut_F2_53[11:0] , REGofMAX1DataOut_F2_54[33:14] } <= AXIinput ; end 
58  + 153 : begin {REGofMAX1DataOut_F2_54[13:0] , REGofMAX1DataOut_F2_55[33:16] } <= AXIinput ; end 
59  + 153 : begin {REGofMAX1DataOut_F2_55[15:0] , REGofMAX1DataOut_F2_56[33:18] } <= AXIinput ; end 
60  + 153 : begin {REGofMAX1DataOut_F2_56[17:0] , REGofMAX1DataOut_F2_57[33:20] } <= AXIinput ; end 
61  + 153 : begin {REGofMAX1DataOut_F2_57[19:0] , REGofMAX1DataOut_F2_58[33:22] } <= AXIinput ; end 
62  + 153 : begin {REGofMAX1DataOut_F2_58[21:0] , REGofMAX1DataOut_F2_59[33:24] } <= AXIinput ; end 
63  + 153 : begin {REGofMAX1DataOut_F2_59[23:0] , REGofMAX1DataOut_F2_60[33:26] } <= AXIinput ; end  
64  + 153 : begin {REGofMAX1DataOut_F2_60[25:0] , REGofMAX1DataOut_F2_61[33:28] } <= AXIinput ; end  
65  + 153 : begin {REGofMAX1DataOut_F2_61[27:0] , REGofMAX1DataOut_F2_62[33:30] } <= AXIinput ; end 
66 + 153 : begin {REGofMAX1DataOut_F2_62[29:0] , REGofMAX1DataOut_F2_63[33:32] } <= AXIinput ; end 
67  + 153 : begin {REGofMAX1DataOut_F2_63[31:0] } <= AXIinput ; end 
68  + 153 : begin {REGofMAX1DataOut_F2_64[33:2] } <= AXIinput ; end 
69  + 153 : begin {REGofMAX1DataOut_F2_64[1:0], REGofMAX1DataOut_F2_65[33:4] } <= AXIinput ; end 
70  + 153 : begin {REGofMAX1DataOut_F2_65[3:0] , REGofMAX1DataOut_F2_66[33:6]  } <= AXIinput ; end  
71  + 153 : begin {REGofMAX1DataOut_F2_66[5:0] , REGofMAX1DataOut_F2_67[33:8]  } <= AXIinput ; end 
72  + 153 : begin {REGofMAX1DataOut_F2_67[7:0] , REGofMAX1DataOut_F2_68[33:10]  } <= AXIinput ; end 
73  + 153 : begin {REGofMAX1DataOut_F2_68[9:0] , REGofMAX1DataOut_F2_69[33:12]  } <= AXIinput ; end 
74  + 153 : begin {REGofMAX1DataOut_F2_69[11:0] , REGofMAX1DataOut_F2_70[33:14] } <= AXIinput ; end 
75  + 153 : begin {REGofMAX1DataOut_F2_70[13:0] , REGofMAX1DataOut_F2_71[33:16] } <= AXIinput ; end 
76  + 153 : begin {REGofMAX1DataOut_F2_71[15:0] , REGofMAX1DataOut_F2_72[33:18] } <= AXIinput ; end  
77  + 153 : begin {REGofMAX1DataOut_F2_72[17:0] , REGofMAX1DataOut_F2_73[33:20] } <= AXIinput ; end 
78  + 153 : begin {REGofMAX1DataOut_F2_73[19:0] , REGofMAX1DataOut_F2_74[33:22] } <= AXIinput ; end 
79  + 153 : begin {REGofMAX1DataOut_F2_74[21:0] , REGofMAX1DataOut_F2_75[33:24] } <= AXIinput ; end 
80  + 153 : begin {REGofMAX1DataOut_F2_75[23:0] , REGofMAX1DataOut_F2_76[33:26] } <= AXIinput ; end 
81  + 153 : begin {REGofMAX1DataOut_F2_76[25:0] , REGofMAX1DataOut_F2_77[33:28] } <= AXIinput ; end 
82  + 153 : begin {REGofMAX1DataOut_F2_77[27:0] , REGofMAX1DataOut_F2_78[33:30] } <= AXIinput ; end 
83  + 153 : begin {REGofMAX1DataOut_F2_78[29:0] , REGofMAX1DataOut_F2_79[33:32] } <= AXIinput ; end 
84  + 153 : begin {REGofMAX1DataOut_F2_79[31:0] } <= AXIinput ; end 
85  + 153 : begin {REGofMAX1DataOut_F2_80[33:2] } <= AXIinput ; end 
86  + 153 : begin {REGofMAX1DataOut_F2_80[1:0], REGofMAX1DataOut_F2_81[33:4] } <= AXIinput ; end 
87  + 153 : begin {REGofMAX1DataOut_F2_81[3:0] , REGofMAX1DataOut_F2_82[33:6]  } <= AXIinput ; end 
88  + 153 : begin {REGofMAX1DataOut_F2_82[5:0] , REGofMAX1DataOut_F2_83[33:8]  } <= AXIinput ; end 
89  + 153 : begin {REGofMAX1DataOut_F2_83[7:0] , REGofMAX1DataOut_F2_84[33:10]  } <= AXIinput ; end 
90  + 153 : begin {REGofMAX1DataOut_F2_84[9:0] , REGofMAX1DataOut_F2_85[33:12]  } <= AXIinput ; end 
91  + 153 : begin {REGofMAX1DataOut_F2_85[11:0] , REGofMAX1DataOut_F2_86[33:14] } <= AXIinput ; end  
92  + 153 : begin {REGofMAX1DataOut_F2_86[13:0] , REGofMAX1DataOut_F2_87[33:16] } <= AXIinput ; end 
93  + 153 : begin {REGofMAX1DataOut_F2_87[15:0] , REGofMAX1DataOut_F2_88[33:18] } <= AXIinput ; end 
94  + 153 : begin {REGofMAX1DataOut_F2_88[17:0] , REGofMAX1DataOut_F2_89[33:20] } <= AXIinput ; end 
95  + 153 : begin {REGofMAX1DataOut_F2_89[19:0] , REGofMAX1DataOut_F2_90[33:22] } <= AXIinput ; end 
96  + 153 : begin {REGofMAX1DataOut_F2_90[21:0] , REGofMAX1DataOut_F2_91[33:24] } <= AXIinput ; end 
97  + 153 : begin {REGofMAX1DataOut_F2_91[23:0] , REGofMAX1DataOut_F2_92[33:26] } <= AXIinput ; end 
98  + 153 : begin {REGofMAX1DataOut_F2_92[25:0] , REGofMAX1DataOut_F2_93[33:28] } <= AXIinput ; end 
99  + 153 : begin {REGofMAX1DataOut_F2_93[27:0] , REGofMAX1DataOut_F2_94[33:30] } <= AXIinput ; end 
100  + 153 : begin {REGofMAX1DataOut_F2_94[29:0] , REGofMAX1DataOut_F2_95[33:32] } <= AXIinput ; end 
101  + 153 : begin {REGofMAX1DataOut_F2_95[31:0] } <= AXIinput ; end 
102  + 153 : begin {REGofMAX1DataOut_F2_96[33:2] } <= AXIinput ; end 
103  + 153 : begin {REGofMAX1DataOut_F2_96[1:0], REGofMAX1DataOut_F2_97[33:4] } <= AXIinput ; end 
104  + 153 : begin {REGofMAX1DataOut_F2_97[3:0] , REGofMAX1DataOut_F2_98[33:6]  } <= AXIinput ; end 
105  + 153 : begin {REGofMAX1DataOut_F2_98[5:0] , REGofMAX1DataOut_F2_99[33:8]  } <= AXIinput ; end  
106  + 153 : begin {REGofMAX1DataOut_F2_99[7:0] , REGofMAX1DataOut_F2_100[33:10]  } <= AXIinput ; end 
107  + 153 : begin {REGofMAX1DataOut_F2_100[9:0] , REGofMAX1DataOut_F2_101[33:12]  } <= AXIinput ; end 
108  + 153 : begin {REGofMAX1DataOut_F2_101[11:0] , REGofMAX1DataOut_F2_102[33:14] } <= AXIinput ; end  
109  + 153 : begin {REGofMAX1DataOut_F2_102[13:0] , REGofMAX1DataOut_F2_103[33:16] } <= AXIinput ; end 
110  + 153 : begin {REGofMAX1DataOut_F2_103[15:0] , REGofMAX1DataOut_F2_104[33:18] } <= AXIinput ; end 
111  + 153 : begin {REGofMAX1DataOut_F2_104[17:0] , REGofMAX1DataOut_F2_105[33:20] } <= AXIinput ; end 
112  + 153 : begin {REGofMAX1DataOut_F2_105[19:0] , REGofMAX1DataOut_F2_106[33:22] } <= AXIinput ; end 
113  + 153 : begin {REGofMAX1DataOut_F2_106[21:0] , REGofMAX1DataOut_F2_107[33:24] } <= AXIinput ; end 
114  + 153 : begin {REGofMAX1DataOut_F2_107[23:0] , REGofMAX1DataOut_F2_108[33:26] } <= AXIinput ; end 
115  + 153 : begin {REGofMAX1DataOut_F2_108[25:0] , REGofMAX1DataOut_F2_109[33:28] } <= AXIinput ; end 
116  + 153 : begin {REGofMAX1DataOut_F2_109[27:0] , REGofMAX1DataOut_F2_110[33:30] } <= AXIinput ; end 
117  + 153 : begin {REGofMAX1DataOut_F2_110[29:0] , REGofMAX1DataOut_F2_111[33:32] } <= AXIinput ; end 
118  + 153 : begin {REGofMAX1DataOut_F2_111[31:0] } <= AXIinput ; end 
119  + 153 : begin {REGofMAX1DataOut_F2_112[33:2] } <= AXIinput ; end 
120  + 153 : begin {REGofMAX1DataOut_F2_112[1:0], REGofMAX1DataOut_F2_113[33:4] } <= AXIinput ; end 
121  + 153 : begin {REGofMAX1DataOut_F2_113[3:0] , REGofMAX1DataOut_F2_114[33:6]  } <= AXIinput ; end 
122  + 153 : begin {REGofMAX1DataOut_F2_114[5:0] , REGofMAX1DataOut_F2_115[33:8]  } <= AXIinput ; end 
123  + 153 : begin {REGofMAX1DataOut_F2_115[7:0] , REGofMAX1DataOut_F2_116[33:10]  } <= AXIinput ; end 
124  + 153 : begin {REGofMAX1DataOut_F2_116[9:0] , REGofMAX1DataOut_F2_117[33:12]  } <= AXIinput ; end 
125  + 153 : begin {REGofMAX1DataOut_F2_117[11:0] , REGofMAX1DataOut_F2_118[33:14] } <= AXIinput ; end 
126  + 153 : begin {REGofMAX1DataOut_F2_118[13:0] , REGofMAX1DataOut_F2_119[33:16] } <= AXIinput ; end 
127  + 153 : begin {REGofMAX1DataOut_F2_119[15:0] , REGofMAX1DataOut_F2_120[33:18] } <= AXIinput ; end 
128  + 153 : begin {REGofMAX1DataOut_F2_120[17:0] , REGofMAX1DataOut_F2_121[33:20] } <= AXIinput ; end 
129  + 153 : begin {REGofMAX1DataOut_F2_121[19:0] , REGofMAX1DataOut_F2_122[33:22] } <= AXIinput ; end 
130  + 153 : begin {REGofMAX1DataOut_F2_122[21:0] , REGofMAX1DataOut_F2_123[33:24] } <= AXIinput ; end 
131  + 153 : begin {REGofMAX1DataOut_F2_123[23:0] , REGofMAX1DataOut_F2_124[33:26] } <= AXIinput ; end 
132  + 153 : begin {REGofMAX1DataOut_F2_124[25:0] , REGofMAX1DataOut_F2_125[33:28] } <= AXIinput ; end 
133  + 153 : begin {REGofMAX1DataOut_F2_125[27:0] , REGofMAX1DataOut_F2_126[33:30] } <= AXIinput ; end 
134  + 153 : begin {REGofMAX1DataOut_F2_126[29:0] , REGofMAX1DataOut_F2_127[33:32] } <= AXIinput ; end 
135  + 153 : begin {REGofMAX1DataOut_F2_127[31:0] } <= AXIinput ; end 
136  + 153 : begin {REGofMAX1DataOut_F2_128[33:2] } <= AXIinput ; end 
137  + 153 : begin {REGofMAX1DataOut_F2_128[1:0], REGofMAX1DataOut_F2_129[33:4] } <= AXIinput ; end 
138  + 153 : begin {REGofMAX1DataOut_F2_129[3:0] , REGofMAX1DataOut_F2_130[33:6]  } <= AXIinput ; end 
139  + 153 : begin {REGofMAX1DataOut_F2_130[5:0] , REGofMAX1DataOut_F2_131[33:8]  } <= AXIinput ; end 
140  + 153 : begin {REGofMAX1DataOut_F2_131[7:0] , REGofMAX1DataOut_F2_132[33:10]  } <= AXIinput ; end 
141  + 153 : begin {REGofMAX1DataOut_F2_132[9:0] , REGofMAX1DataOut_F2_133[33:12]  } <= AXIinput ; end 
142  + 153 : begin {REGofMAX1DataOut_F2_133[11:0] , REGofMAX1DataOut_F2_134[33:14] } <= AXIinput ; end 
143  + 153 : begin {REGofMAX1DataOut_F2_134[13:0] , REGofMAX1DataOut_F2_135[33:16] } <= AXIinput ; end 
144  + 153 : begin {REGofMAX1DataOut_F2_135[15:0] , REGofMAX1DataOut_F2_136[33:18] } <= AXIinput ; end 
145  + 153 : begin {REGofMAX1DataOut_F2_136[17:0] , REGofMAX1DataOut_F2_137[33:20] } <= AXIinput ; end 
146  + 153 : begin {REGofMAX1DataOut_F2_137[19:0] , REGofMAX1DataOut_F2_138[33:22] } <= AXIinput ; end 
147  + 153 : begin {REGofMAX1DataOut_F2_138[21:0] , REGofMAX1DataOut_F2_139[33:24] } <= AXIinput ; end 
148  + 153 : begin {REGofMAX1DataOut_F2_139[23:0] , REGofMAX1DataOut_F2_140[33:26] } <= AXIinput ; end 
149  + 153 : begin {REGofMAX1DataOut_F2_140[25:0] , REGofMAX1DataOut_F2_141[33:28] } <= AXIinput ; end 
150  + 153 : begin {REGofMAX1DataOut_F2_141[27:0] , REGofMAX1DataOut_F2_142[33:30] } <= AXIinput ; end 
151  + 153 : begin {REGofMAX1DataOut_F2_142[29:0] , REGofMAX1DataOut_F2_143[33:32] } <= AXIinput ; end 
152  + 153 : begin {REGofMAX1DataOut_F2_143[31:0] } <= AXIinput ; end 


0  + 306 : begin {REGofMAX1DataOut_F3_0[33:2] } <= AXIinput ; end 
1  + 306 : begin {REGofMAX1DataOut_F3_0[1:0] , REGofMAX1DataOut_F3_1[33:4] } <= AXIinput ; end 
2  + 306 : begin {REGofMAX1DataOut_F3_1[3:0] , REGofMAX1DataOut_F3_2[33:6]  } <= AXIinput ; end 
3  + 306 : begin {REGofMAX1DataOut_F3_2[5:0] , REGofMAX1DataOut_F3_3[33:8]  } <= AXIinput ; end 
4  + 306 : begin {REGofMAX1DataOut_F3_3[7:0] , REGofMAX1DataOut_F3_4[33:10]  } <= AXIinput ; end 
5  + 306 : begin {REGofMAX1DataOut_F3_4[9:0] , REGofMAX1DataOut_F3_5[33:12]  } <= AXIinput ; end 
6  + 306 : begin {REGofMAX1DataOut_F3_5[11:0] , REGofMAX1DataOut_F3_6[33:14] } <= AXIinput ; end 
7  + 306 : begin {REGofMAX1DataOut_F3_6[13:0] , REGofMAX1DataOut_F3_7[33:16] } <= AXIinput ; end 
8  + 306 : begin {REGofMAX1DataOut_F3_7[15:0] , REGofMAX1DataOut_F3_8[33:18] } <= AXIinput ; end 
9  + 306 : begin {REGofMAX1DataOut_F3_8[17:0] , REGofMAX1DataOut_F3_9[33:20] } <= AXIinput ; end 
10  + 306 : begin {REGofMAX1DataOut_F3_9[19:0] , REGofMAX1DataOut_F3_10[33:22] } <= AXIinput ; end 
11  + 306 : begin {REGofMAX1DataOut_F3_10[21:0] , REGofMAX1DataOut_F3_11[33:24] } <= AXIinput ; end  
12  + 306 : begin {REGofMAX1DataOut_F3_11[23:0] , REGofMAX1DataOut_F3_12[33:26] } <= AXIinput ; end 
13  + 306 : begin {REGofMAX1DataOut_F3_12[25:0] , REGofMAX1DataOut_F3_13[33:28] } <= AXIinput ; end 
14  + 306 : begin {REGofMAX1DataOut_F3_13[27:0] , REGofMAX1DataOut_F3_14[33:30] } <= AXIinput ; end 
15  + 306 : begin {REGofMAX1DataOut_F3_14[29:0] , REGofMAX1DataOut_F3_15[33:32] } <= AXIinput ; end 
16  + 306 : begin {REGofMAX1DataOut_F3_15[31:0] } <= AXIinput ; end 
17  + 306 : begin {REGofMAX1DataOut_F3_16[33:2] } <= AXIinput ; end 
18  + 306 : begin {REGofMAX1DataOut_F3_16[1:0], REGofMAX1DataOut_F3_17[33:4] } <= AXIinput ; end 
19  + 306 : begin {REGofMAX1DataOut_F3_17[3:0] , REGofMAX1DataOut_F3_18[33:6]  } <= AXIinput ; end 
20  + 306 : begin {REGofMAX1DataOut_F3_18[5:0] , REGofMAX1DataOut_F3_19[33:8]  } <= AXIinput ; end 
21  + 306 : begin {REGofMAX1DataOut_F3_19[7:0] , REGofMAX1DataOut_F3_20[33:10]  } <= AXIinput ; end 
22  + 306 : begin {REGofMAX1DataOut_F3_20[9:0] , REGofMAX1DataOut_F3_21[33:12]  } <= AXIinput ; end 
23  + 306 : begin {REGofMAX1DataOut_F3_21[11:0] , REGofMAX1DataOut_F3_22[33:14] } <= AXIinput ; end 
24  + 306 : begin {REGofMAX1DataOut_F3_22[13:0] , REGofMAX1DataOut_F3_23[33:16] } <= AXIinput ; end 
25  + 306 : begin {REGofMAX1DataOut_F3_23[15:0] , REGofMAX1DataOut_F3_24[33:18] } <= AXIinput ; end 
26  + 306 : begin {REGofMAX1DataOut_F3_24[17:0] , REGofMAX1DataOut_F3_25[33:20] } <= AXIinput ; end 
27  + 306 : begin {REGofMAX1DataOut_F3_25[19:0] , REGofMAX1DataOut_F3_26[33:22] } <= AXIinput ; end 
28  + 306 : begin {REGofMAX1DataOut_F3_26[21:0] , REGofMAX1DataOut_F3_27[33:24] } <= AXIinput ; end  
29  + 306 : begin {REGofMAX1DataOut_F3_27[23:0] , REGofMAX1DataOut_F3_28[33:26] } <= AXIinput ; end 
30  + 306 : begin {REGofMAX1DataOut_F3_28[25:0] , REGofMAX1DataOut_F3_29[33:28] } <= AXIinput ; end 
31  + 306 : begin {REGofMAX1DataOut_F3_29[27:0] , REGofMAX1DataOut_F3_30[33:30] } <= AXIinput ; end 
32  + 306 : begin {REGofMAX1DataOut_F3_30[29:0] , REGofMAX1DataOut_F3_31[33:32] } <= AXIinput ; end 
33  + 306 : begin {REGofMAX1DataOut_F3_31[31:0] } <= AXIinput ; end 
34  + 306 : begin {REGofMAX1DataOut_F3_32[33:2] } <= AXIinput ; end 
35  + 306 : begin {REGofMAX1DataOut_F3_32[1:0], REGofMAX1DataOut_F3_33[33:4] } <= AXIinput ; end 
36  + 306 : begin {REGofMAX1DataOut_F3_33[3:0] , REGofMAX1DataOut_F3_34[33:6]  } <= AXIinput ; end 
37  + 306 : begin {REGofMAX1DataOut_F3_34[5:0] , REGofMAX1DataOut_F3_35[33:8]  } <= AXIinput ; end 
38  + 306 : begin {REGofMAX1DataOut_F3_35[7:0] , REGofMAX1DataOut_F3_36[33:10]  } <= AXIinput ; end 
39  + 306 : begin {REGofMAX1DataOut_F3_36[9:0] , REGofMAX1DataOut_F3_37[33:12]  } <= AXIinput ; end 
40  + 306 : begin {REGofMAX1DataOut_F3_37[11:0] , REGofMAX1DataOut_F3_38[33:14] } <= AXIinput ; end  
41  + 306 : begin {REGofMAX1DataOut_F3_38[13:0] , REGofMAX1DataOut_F3_39[33:16] } <= AXIinput ; end 
42  + 306 : begin {REGofMAX1DataOut_F3_39[15:0] , REGofMAX1DataOut_F3_40[33:18] } <= AXIinput ; end 
43  + 306 : begin {REGofMAX1DataOut_F3_40[17:0] , REGofMAX1DataOut_F3_41[33:20] } <= AXIinput ; end 
44  + 306 : begin {REGofMAX1DataOut_F3_41[19:0] , REGofMAX1DataOut_F3_42[33:22] } <= AXIinput ; end  
45  + 306 : begin {REGofMAX1DataOut_F3_42[21:0] , REGofMAX1DataOut_F3_43[33:24] } <= AXIinput ; end 
46  + 306 : begin {REGofMAX1DataOut_F3_43[23:0] , REGofMAX1DataOut_F3_44[33:26] } <= AXIinput ; end 
47  + 306 : begin {REGofMAX1DataOut_F3_44[25:0] , REGofMAX1DataOut_F3_45[33:28] } <= AXIinput ; end  
48  + 306 : begin {REGofMAX1DataOut_F3_45[27:0] , REGofMAX1DataOut_F3_46[33:30] } <= AXIinput ; end 
49  + 306 : begin {REGofMAX1DataOut_F3_46[29:0] , REGofMAX1DataOut_F3_47[33:32] } <= AXIinput ; end 
50  + 306 : begin {REGofMAX1DataOut_F3_47[31:0] } <= AXIinput ; end
51  + 306 : begin {REGofMAX1DataOut_F3_48[33:2] } <= AXIinput ; end 
52  + 306 : begin {REGofMAX1DataOut_F3_48[1:0], REGofMAX1DataOut_F3_49[33:4] } <= AXIinput ; end 
53  + 306 : begin {REGofMAX1DataOut_F3_49[3:0] , REGofMAX1DataOut_F3_50[33:6]  } <= AXIinput ; end 
54  + 306 : begin {REGofMAX1DataOut_F3_50[5:0] , REGofMAX1DataOut_F3_51[33:8]  } <= AXIinput ; end 
55  + 306 : begin {REGofMAX1DataOut_F3_51[7:0] , REGofMAX1DataOut_F3_52[33:10]  } <= AXIinput ; end 
56  + 306 : begin {REGofMAX1DataOut_F3_52[9:0] , REGofMAX1DataOut_F3_53[33:12]  } <= AXIinput ; end 
57  + 306 : begin {REGofMAX1DataOut_F3_53[11:0] , REGofMAX1DataOut_F3_54[33:14] } <= AXIinput ; end 
58  + 306 : begin {REGofMAX1DataOut_F3_54[13:0] , REGofMAX1DataOut_F3_55[33:16] } <= AXIinput ; end 
59  + 306 : begin {REGofMAX1DataOut_F3_55[15:0] , REGofMAX1DataOut_F3_56[33:18] } <= AXIinput ; end 
60  + 306 : begin {REGofMAX1DataOut_F3_56[17:0] , REGofMAX1DataOut_F3_57[33:20] } <= AXIinput ; end 
61  + 306 : begin {REGofMAX1DataOut_F3_57[19:0] , REGofMAX1DataOut_F3_58[33:22] } <= AXIinput ; end 
62  + 306 : begin {REGofMAX1DataOut_F3_58[21:0] , REGofMAX1DataOut_F3_59[33:24] } <= AXIinput ; end 
63  + 306 : begin {REGofMAX1DataOut_F3_59[23:0] , REGofMAX1DataOut_F3_60[33:26] } <= AXIinput ; end  
64  + 306 : begin {REGofMAX1DataOut_F3_60[25:0] , REGofMAX1DataOut_F3_61[33:28] } <= AXIinput ; end  
65  + 306 : begin {REGofMAX1DataOut_F3_61[27:0] , REGofMAX1DataOut_F3_62[33:30] } <= AXIinput ; end 
66 + 306 : begin {REGofMAX1DataOut_F3_62[29:0] , REGofMAX1DataOut_F3_63[33:32] } <= AXIinput ; end 
67  + 306 : begin {REGofMAX1DataOut_F3_63[31:0] } <= AXIinput ; end 
68  + 306 : begin {REGofMAX1DataOut_F3_64[33:2] } <= AXIinput ; end 
69  + 306 : begin {REGofMAX1DataOut_F3_64[1:0], REGofMAX1DataOut_F3_65[33:4] } <= AXIinput ; end 
70  + 306 : begin {REGofMAX1DataOut_F3_65[3:0] , REGofMAX1DataOut_F3_66[33:6]  } <= AXIinput ; end  
71  + 306 : begin {REGofMAX1DataOut_F3_66[5:0] , REGofMAX1DataOut_F3_67[33:8]  } <= AXIinput ; end 
72  + 306 : begin {REGofMAX1DataOut_F3_67[7:0] , REGofMAX1DataOut_F3_68[33:10]  } <= AXIinput ; end 
73  + 306 : begin {REGofMAX1DataOut_F3_68[9:0] , REGofMAX1DataOut_F3_69[33:12]  } <= AXIinput ; end 
74  + 306 : begin {REGofMAX1DataOut_F3_69[11:0] , REGofMAX1DataOut_F3_70[33:14] } <= AXIinput ; end 
75  + 306 : begin {REGofMAX1DataOut_F3_70[13:0] , REGofMAX1DataOut_F3_71[33:16] } <= AXIinput ; end 
76  + 306 : begin {REGofMAX1DataOut_F3_71[15:0] , REGofMAX1DataOut_F3_72[33:18] } <= AXIinput ; end  
77  + 306 : begin {REGofMAX1DataOut_F3_72[17:0] , REGofMAX1DataOut_F3_73[33:20] } <= AXIinput ; end 
78  + 306 : begin {REGofMAX1DataOut_F3_73[19:0] , REGofMAX1DataOut_F3_74[33:22] } <= AXIinput ; end 
79  + 306 : begin {REGofMAX1DataOut_F3_74[21:0] , REGofMAX1DataOut_F3_75[33:24] } <= AXIinput ; end 
80  + 306 : begin {REGofMAX1DataOut_F3_75[23:0] , REGofMAX1DataOut_F3_76[33:26] } <= AXIinput ; end 
81  + 306 : begin {REGofMAX1DataOut_F3_76[25:0] , REGofMAX1DataOut_F3_77[33:28] } <= AXIinput ; end 
82  + 306 : begin {REGofMAX1DataOut_F3_77[27:0] , REGofMAX1DataOut_F3_78[33:30] } <= AXIinput ; end 
83  + 306 : begin {REGofMAX1DataOut_F3_78[29:0] , REGofMAX1DataOut_F3_79[33:32] } <= AXIinput ; end 
84  + 306 : begin {REGofMAX1DataOut_F3_79[31:0] } <= AXIinput ; end 
85  + 306 : begin {REGofMAX1DataOut_F3_80[33:2] } <= AXIinput ; end 
86  + 306 : begin {REGofMAX1DataOut_F3_80[1:0], REGofMAX1DataOut_F3_81[33:4] } <= AXIinput ; end 
87  + 306 : begin {REGofMAX1DataOut_F3_81[3:0] , REGofMAX1DataOut_F3_82[33:6]  } <= AXIinput ; end 
88  + 306 : begin {REGofMAX1DataOut_F3_82[5:0] , REGofMAX1DataOut_F3_83[33:8]  } <= AXIinput ; end 
89  + 306 : begin {REGofMAX1DataOut_F3_83[7:0] , REGofMAX1DataOut_F3_84[33:10]  } <= AXIinput ; end 
90  + 306 : begin {REGofMAX1DataOut_F3_84[9:0] , REGofMAX1DataOut_F3_85[33:12]  } <= AXIinput ; end 
91  + 306 : begin {REGofMAX1DataOut_F3_85[11:0] , REGofMAX1DataOut_F3_86[33:14] } <= AXIinput ; end  
92  + 306 : begin {REGofMAX1DataOut_F3_86[13:0] , REGofMAX1DataOut_F3_87[33:16] } <= AXIinput ; end 
93  + 306 : begin {REGofMAX1DataOut_F3_87[15:0] , REGofMAX1DataOut_F3_88[33:18] } <= AXIinput ; end 
94  + 306 : begin {REGofMAX1DataOut_F3_88[17:0] , REGofMAX1DataOut_F3_89[33:20] } <= AXIinput ; end 
95  + 306 : begin {REGofMAX1DataOut_F3_89[19:0] , REGofMAX1DataOut_F3_90[33:22] } <= AXIinput ; end 
96  + 306 : begin {REGofMAX1DataOut_F3_90[21:0] , REGofMAX1DataOut_F3_91[33:24] } <= AXIinput ; end 
97  + 306 : begin {REGofMAX1DataOut_F3_91[23:0] , REGofMAX1DataOut_F3_92[33:26] } <= AXIinput ; end 
98  + 306 : begin {REGofMAX1DataOut_F3_92[25:0] , REGofMAX1DataOut_F3_93[33:28] } <= AXIinput ; end 
99  + 306 : begin {REGofMAX1DataOut_F3_93[27:0] , REGofMAX1DataOut_F3_94[33:30] } <= AXIinput ; end 
100  + 306 : begin {REGofMAX1DataOut_F3_94[29:0] , REGofMAX1DataOut_F3_95[33:32] } <= AXIinput ; end 
101  + 306 : begin {REGofMAX1DataOut_F3_95[31:0] } <= AXIinput ; end 
102  + 306 : begin {REGofMAX1DataOut_F3_96[33:2] } <= AXIinput ; end 
103  + 306 : begin {REGofMAX1DataOut_F3_96[1:0], REGofMAX1DataOut_F3_97[33:4] } <= AXIinput ; end 
104  + 306 : begin {REGofMAX1DataOut_F3_97[3:0] , REGofMAX1DataOut_F3_98[33:6]  } <= AXIinput ; end 
105  + 306 : begin {REGofMAX1DataOut_F3_98[5:0] , REGofMAX1DataOut_F3_99[33:8]  } <= AXIinput ; end  
106  + 306 : begin {REGofMAX1DataOut_F3_99[7:0] , REGofMAX1DataOut_F3_100[33:10]  } <= AXIinput ; end 
107  + 306 : begin {REGofMAX1DataOut_F3_100[9:0] , REGofMAX1DataOut_F3_101[33:12]  } <= AXIinput ; end 
108  + 306 : begin {REGofMAX1DataOut_F3_101[11:0] , REGofMAX1DataOut_F3_102[33:14] } <= AXIinput ; end  
109  + 306 : begin {REGofMAX1DataOut_F3_102[13:0] , REGofMAX1DataOut_F3_103[33:16] } <= AXIinput ; end 
110  + 306 : begin {REGofMAX1DataOut_F3_103[15:0] , REGofMAX1DataOut_F3_104[33:18] } <= AXIinput ; end 
111  + 306 : begin {REGofMAX1DataOut_F3_104[17:0] , REGofMAX1DataOut_F3_105[33:20] } <= AXIinput ; end 
112  + 306 : begin {REGofMAX1DataOut_F3_105[19:0] , REGofMAX1DataOut_F3_106[33:22] } <= AXIinput ; end 
113  + 306 : begin {REGofMAX1DataOut_F3_106[21:0] , REGofMAX1DataOut_F3_107[33:24] } <= AXIinput ; end 
114  + 306 : begin {REGofMAX1DataOut_F3_107[23:0] , REGofMAX1DataOut_F3_108[33:26] } <= AXIinput ; end 
115  + 306 : begin {REGofMAX1DataOut_F3_108[25:0] , REGofMAX1DataOut_F3_109[33:28] } <= AXIinput ; end 
116  + 306 : begin {REGofMAX1DataOut_F3_109[27:0] , REGofMAX1DataOut_F3_110[33:30] } <= AXIinput ; end 
117  + 306 : begin {REGofMAX1DataOut_F3_110[29:0] , REGofMAX1DataOut_F3_111[33:32] } <= AXIinput ; end 
118  + 306 : begin {REGofMAX1DataOut_F3_111[31:0] } <= AXIinput ; end 
119  + 306 : begin {REGofMAX1DataOut_F3_112[33:2] } <= AXIinput ; end 
120  + 306 : begin {REGofMAX1DataOut_F3_112[1:0], REGofMAX1DataOut_F3_113[33:4] } <= AXIinput ; end 
121  + 306 : begin {REGofMAX1DataOut_F3_113[3:0] , REGofMAX1DataOut_F3_114[33:6]  } <= AXIinput ; end 
122  + 306 : begin {REGofMAX1DataOut_F3_114[5:0] , REGofMAX1DataOut_F3_115[33:8]  } <= AXIinput ; end 
123  + 306 : begin {REGofMAX1DataOut_F3_115[7:0] , REGofMAX1DataOut_F3_116[33:10]  } <= AXIinput ; end 
124  + 306 : begin {REGofMAX1DataOut_F3_116[9:0] , REGofMAX1DataOut_F3_117[33:12]  } <= AXIinput ; end 
125  + 306 : begin {REGofMAX1DataOut_F3_117[11:0] , REGofMAX1DataOut_F3_118[33:14] } <= AXIinput ; end 
126  + 306 : begin {REGofMAX1DataOut_F3_118[13:0] , REGofMAX1DataOut_F3_119[33:16] } <= AXIinput ; end 
127  + 306 : begin {REGofMAX1DataOut_F3_119[15:0] , REGofMAX1DataOut_F3_120[33:18] } <= AXIinput ; end 
128  + 306 : begin {REGofMAX1DataOut_F3_120[17:0] , REGofMAX1DataOut_F3_121[33:20] } <= AXIinput ; end 
129  + 306 : begin {REGofMAX1DataOut_F3_121[19:0] , REGofMAX1DataOut_F3_122[33:22] } <= AXIinput ; end 
130  + 306 : begin {REGofMAX1DataOut_F3_122[21:0] , REGofMAX1DataOut_F3_123[33:24] } <= AXIinput ; end 
131  + 306 : begin {REGofMAX1DataOut_F3_123[23:0] , REGofMAX1DataOut_F3_124[33:26] } <= AXIinput ; end 
132  + 306 : begin {REGofMAX1DataOut_F3_124[25:0] , REGofMAX1DataOut_F3_125[33:28] } <= AXIinput ; end 
133  + 306 : begin {REGofMAX1DataOut_F3_125[27:0] , REGofMAX1DataOut_F3_126[33:30] } <= AXIinput ; end 
134  + 306 : begin {REGofMAX1DataOut_F3_126[29:0] , REGofMAX1DataOut_F3_127[33:32] } <= AXIinput ; end 
135  + 306 : begin {REGofMAX1DataOut_F3_127[31:0] } <= AXIinput ; end 
136  + 306 : begin {REGofMAX1DataOut_F3_128[33:2] } <= AXIinput ; end 
137  + 306 : begin {REGofMAX1DataOut_F3_128[1:0], REGofMAX1DataOut_F3_129[33:4] } <= AXIinput ; end 
138  + 306 : begin {REGofMAX1DataOut_F3_129[3:0] , REGofMAX1DataOut_F3_130[33:6]  } <= AXIinput ; end 
139  + 306 : begin {REGofMAX1DataOut_F3_130[5:0] , REGofMAX1DataOut_F3_131[33:8]  } <= AXIinput ; end 
140  + 306 : begin {REGofMAX1DataOut_F3_131[7:0] , REGofMAX1DataOut_F3_132[33:10]  } <= AXIinput ; end 
141  + 306 : begin {REGofMAX1DataOut_F3_132[9:0] , REGofMAX1DataOut_F3_133[33:12]  } <= AXIinput ; end 
142  + 306 : begin {REGofMAX1DataOut_F3_133[11:0] , REGofMAX1DataOut_F3_134[33:14] } <= AXIinput ; end 
143  + 306 : begin {REGofMAX1DataOut_F3_134[13:0] , REGofMAX1DataOut_F3_135[33:16] } <= AXIinput ; end 
144  + 306 : begin {REGofMAX1DataOut_F3_135[15:0] , REGofMAX1DataOut_F3_136[33:18] } <= AXIinput ; end 
145  + 306 : begin {REGofMAX1DataOut_F3_136[17:0] , REGofMAX1DataOut_F3_137[33:20] } <= AXIinput ; end 
146  + 306 : begin {REGofMAX1DataOut_F3_137[19:0] , REGofMAX1DataOut_F3_138[33:22] } <= AXIinput ; end 
147  + 306 : begin {REGofMAX1DataOut_F3_138[21:0] , REGofMAX1DataOut_F3_139[33:24] } <= AXIinput ; end 
148  + 306 : begin {REGofMAX1DataOut_F3_139[23:0] , REGofMAX1DataOut_F3_140[33:26] } <= AXIinput ; end 
149  + 306 : begin {REGofMAX1DataOut_F3_140[25:0] , REGofMAX1DataOut_F3_141[33:28] } <= AXIinput ; end 
150  + 306 : begin {REGofMAX1DataOut_F3_141[27:0] , REGofMAX1DataOut_F3_142[33:30] } <= AXIinput ; end 
151  + 306 : begin {REGofMAX1DataOut_F3_142[29:0] , REGofMAX1DataOut_F3_143[33:32] } <= AXIinput ; end 
152  + 306 : begin {REGofMAX1DataOut_F3_143[31:0] } <= AXIinput ; end 


0  + 459 : begin {REGofMAX1DataOut_F4_0[33:2] } <= AXIinput ; end 
1  + 459 : begin {REGofMAX1DataOut_F4_0[1:0] , REGofMAX1DataOut_F4_1[33:4] } <= AXIinput ; end 
2  + 459 : begin {REGofMAX1DataOut_F4_1[3:0] , REGofMAX1DataOut_F4_2[33:6]  } <= AXIinput ; end 
3  + 459 : begin {REGofMAX1DataOut_F4_2[5:0] , REGofMAX1DataOut_F4_3[33:8]  } <= AXIinput ; end 
4  + 459 : begin {REGofMAX1DataOut_F4_3[7:0] , REGofMAX1DataOut_F4_4[33:10]  } <= AXIinput ; end 
5  + 459 : begin {REGofMAX1DataOut_F4_4[9:0] , REGofMAX1DataOut_F4_5[33:12]  } <= AXIinput ; end 
6  + 459 : begin {REGofMAX1DataOut_F4_5[11:0] , REGofMAX1DataOut_F4_6[33:14] } <= AXIinput ; end 
7  + 459 : begin {REGofMAX1DataOut_F4_6[13:0] , REGofMAX1DataOut_F4_7[33:16] } <= AXIinput ; end 
8  + 459 : begin {REGofMAX1DataOut_F4_7[15:0] , REGofMAX1DataOut_F4_8[33:18] } <= AXIinput ; end 
9  + 459 : begin {REGofMAX1DataOut_F4_8[17:0] , REGofMAX1DataOut_F4_9[33:20] } <= AXIinput ; end 
10  + 459 : begin {REGofMAX1DataOut_F4_9[19:0] , REGofMAX1DataOut_F4_10[33:22] } <= AXIinput ; end 
11  + 459 : begin {REGofMAX1DataOut_F4_10[21:0] , REGofMAX1DataOut_F4_11[33:24] } <= AXIinput ; end  
12  + 459 : begin {REGofMAX1DataOut_F4_11[23:0] , REGofMAX1DataOut_F4_12[33:26] } <= AXIinput ; end 
13  + 459 : begin {REGofMAX1DataOut_F4_12[25:0] , REGofMAX1DataOut_F4_13[33:28] } <= AXIinput ; end 
14  + 459 : begin {REGofMAX1DataOut_F4_13[27:0] , REGofMAX1DataOut_F4_14[33:30] } <= AXIinput ; end 
15  + 459 : begin {REGofMAX1DataOut_F4_14[29:0] , REGofMAX1DataOut_F4_15[33:32] } <= AXIinput ; end 
16  + 459 : begin {REGofMAX1DataOut_F4_15[31:0] } <= AXIinput ; end 
17  + 459 : begin {REGofMAX1DataOut_F4_16[33:2] } <= AXIinput ; end 
18  + 459 : begin {REGofMAX1DataOut_F4_16[1:0], REGofMAX1DataOut_F4_17[33:4] } <= AXIinput ; end 
19  + 459 : begin {REGofMAX1DataOut_F4_17[3:0] , REGofMAX1DataOut_F4_18[33:6]  } <= AXIinput ; end 
20  + 459 : begin {REGofMAX1DataOut_F4_18[5:0] , REGofMAX1DataOut_F4_19[33:8]  } <= AXIinput ; end 
21  + 459 : begin {REGofMAX1DataOut_F4_19[7:0] , REGofMAX1DataOut_F4_20[33:10]  } <= AXIinput ; end 
22  + 459 : begin {REGofMAX1DataOut_F4_20[9:0] , REGofMAX1DataOut_F4_21[33:12]  } <= AXIinput ; end 
23  + 459 : begin {REGofMAX1DataOut_F4_21[11:0] , REGofMAX1DataOut_F4_22[33:14] } <= AXIinput ; end 
24  + 459 : begin {REGofMAX1DataOut_F4_22[13:0] , REGofMAX1DataOut_F4_23[33:16] } <= AXIinput ; end 
25  + 459 : begin {REGofMAX1DataOut_F4_23[15:0] , REGofMAX1DataOut_F4_24[33:18] } <= AXIinput ; end 
26  + 459 : begin {REGofMAX1DataOut_F4_24[17:0] , REGofMAX1DataOut_F4_25[33:20] } <= AXIinput ; end 
27  + 459 : begin {REGofMAX1DataOut_F4_25[19:0] , REGofMAX1DataOut_F4_26[33:22] } <= AXIinput ; end 
28  + 459 : begin {REGofMAX1DataOut_F4_26[21:0] , REGofMAX1DataOut_F4_27[33:24] } <= AXIinput ; end  
29  + 459 : begin {REGofMAX1DataOut_F4_27[23:0] , REGofMAX1DataOut_F4_28[33:26] } <= AXIinput ; end 
30  + 459 : begin {REGofMAX1DataOut_F4_28[25:0] , REGofMAX1DataOut_F4_29[33:28] } <= AXIinput ; end 
31  + 459 : begin {REGofMAX1DataOut_F4_29[27:0] , REGofMAX1DataOut_F4_30[33:30] } <= AXIinput ; end 
32  + 459 : begin {REGofMAX1DataOut_F4_30[29:0] , REGofMAX1DataOut_F4_31[33:32] } <= AXIinput ; end 
33  + 459 : begin {REGofMAX1DataOut_F4_31[31:0] } <= AXIinput ; end 
34  + 459 : begin {REGofMAX1DataOut_F4_32[33:2] } <= AXIinput ; end 
35  + 459 : begin {REGofMAX1DataOut_F4_32[1:0], REGofMAX1DataOut_F4_33[33:4] } <= AXIinput ; end 
36  + 459 : begin {REGofMAX1DataOut_F4_33[3:0] , REGofMAX1DataOut_F4_34[33:6]  } <= AXIinput ; end 
37  + 459 : begin {REGofMAX1DataOut_F4_34[5:0] , REGofMAX1DataOut_F4_35[33:8]  } <= AXIinput ; end 
38  + 459 : begin {REGofMAX1DataOut_F4_35[7:0] , REGofMAX1DataOut_F4_36[33:10]  } <= AXIinput ; end 
39  + 459 : begin {REGofMAX1DataOut_F4_36[9:0] , REGofMAX1DataOut_F4_37[33:12]  } <= AXIinput ; end 
40  + 459 : begin {REGofMAX1DataOut_F4_37[11:0] , REGofMAX1DataOut_F4_38[33:14] } <= AXIinput ; end  
41  + 459 : begin {REGofMAX1DataOut_F4_38[13:0] , REGofMAX1DataOut_F4_39[33:16] } <= AXIinput ; end 
42  + 459 : begin {REGofMAX1DataOut_F4_39[15:0] , REGofMAX1DataOut_F4_40[33:18] } <= AXIinput ; end 
43  + 459 : begin {REGofMAX1DataOut_F4_40[17:0] , REGofMAX1DataOut_F4_41[33:20] } <= AXIinput ; end 
44  + 459 : begin {REGofMAX1DataOut_F4_41[19:0] , REGofMAX1DataOut_F4_42[33:22] } <= AXIinput ; end  
45  + 459 : begin {REGofMAX1DataOut_F4_42[21:0] , REGofMAX1DataOut_F4_43[33:24] } <= AXIinput ; end 
46  + 459 : begin {REGofMAX1DataOut_F4_43[23:0] , REGofMAX1DataOut_F4_44[33:26] } <= AXIinput ; end 
47  + 459 : begin {REGofMAX1DataOut_F4_44[25:0] , REGofMAX1DataOut_F4_45[33:28] } <= AXIinput ; end  
48  + 459 : begin {REGofMAX1DataOut_F4_45[27:0] , REGofMAX1DataOut_F4_46[33:30] } <= AXIinput ; end 
49  + 459 : begin {REGofMAX1DataOut_F4_46[29:0] , REGofMAX1DataOut_F4_47[33:32] } <= AXIinput ; end 
50  + 459 : begin {REGofMAX1DataOut_F4_47[31:0] } <= AXIinput ; end
51  + 459 : begin {REGofMAX1DataOut_F4_48[33:2] } <= AXIinput ; end 
52  + 459 : begin {REGofMAX1DataOut_F4_48[1:0], REGofMAX1DataOut_F4_49[33:4] } <= AXIinput ; end 
53  + 459 : begin {REGofMAX1DataOut_F4_49[3:0] , REGofMAX1DataOut_F4_50[33:6]  } <= AXIinput ; end 
54  + 459 : begin {REGofMAX1DataOut_F4_50[5:0] , REGofMAX1DataOut_F4_51[33:8]  } <= AXIinput ; end 
55  + 459 : begin {REGofMAX1DataOut_F4_51[7:0] , REGofMAX1DataOut_F4_52[33:10]  } <= AXIinput ; end 
56  + 459 : begin {REGofMAX1DataOut_F4_52[9:0] , REGofMAX1DataOut_F4_53[33:12]  } <= AXIinput ; end 
57  + 459 : begin {REGofMAX1DataOut_F4_53[11:0] , REGofMAX1DataOut_F4_54[33:14] } <= AXIinput ; end 
58  + 459 : begin {REGofMAX1DataOut_F4_54[13:0] , REGofMAX1DataOut_F4_55[33:16] } <= AXIinput ; end 
59  + 459 : begin {REGofMAX1DataOut_F4_55[15:0] , REGofMAX1DataOut_F4_56[33:18] } <= AXIinput ; end 
60  + 459 : begin {REGofMAX1DataOut_F4_56[17:0] , REGofMAX1DataOut_F4_57[33:20] } <= AXIinput ; end 
61  + 459 : begin {REGofMAX1DataOut_F4_57[19:0] , REGofMAX1DataOut_F4_58[33:22] } <= AXIinput ; end 
62  + 459 : begin {REGofMAX1DataOut_F4_58[21:0] , REGofMAX1DataOut_F4_59[33:24] } <= AXIinput ; end 
63  + 459 : begin {REGofMAX1DataOut_F4_59[23:0] , REGofMAX1DataOut_F4_60[33:26] } <= AXIinput ; end  
64  + 459 : begin {REGofMAX1DataOut_F4_60[25:0] , REGofMAX1DataOut_F4_61[33:28] } <= AXIinput ; end  
65  + 459 : begin {REGofMAX1DataOut_F4_61[27:0] , REGofMAX1DataOut_F4_62[33:30] } <= AXIinput ; end 
66 + 459 : begin {REGofMAX1DataOut_F4_62[29:0] , REGofMAX1DataOut_F4_63[33:32] } <= AXIinput ; end 
67  + 459 : begin {REGofMAX1DataOut_F4_63[31:0] } <= AXIinput ; end 
68  + 459 : begin {REGofMAX1DataOut_F4_64[33:2] } <= AXIinput ; end 
69  + 459 : begin {REGofMAX1DataOut_F4_64[1:0], REGofMAX1DataOut_F4_65[33:4] } <= AXIinput ; end 
70  + 459 : begin {REGofMAX1DataOut_F4_65[3:0] , REGofMAX1DataOut_F4_66[33:6]  } <= AXIinput ; end  
71  + 459 : begin {REGofMAX1DataOut_F4_66[5:0] , REGofMAX1DataOut_F4_67[33:8]  } <= AXIinput ; end 
72  + 459 : begin {REGofMAX1DataOut_F4_67[7:0] , REGofMAX1DataOut_F4_68[33:10]  } <= AXIinput ; end 
73  + 459 : begin {REGofMAX1DataOut_F4_68[9:0] , REGofMAX1DataOut_F4_69[33:12]  } <= AXIinput ; end 
74  + 459 : begin {REGofMAX1DataOut_F4_69[11:0] , REGofMAX1DataOut_F4_70[33:14] } <= AXIinput ; end 
75  + 459 : begin {REGofMAX1DataOut_F4_70[13:0] , REGofMAX1DataOut_F4_71[33:16] } <= AXIinput ; end 
76  + 459 : begin {REGofMAX1DataOut_F4_71[15:0] , REGofMAX1DataOut_F4_72[33:18] } <= AXIinput ; end  
77  + 459 : begin {REGofMAX1DataOut_F4_72[17:0] , REGofMAX1DataOut_F4_73[33:20] } <= AXIinput ; end 
78  + 459 : begin {REGofMAX1DataOut_F4_73[19:0] , REGofMAX1DataOut_F4_74[33:22] } <= AXIinput ; end 
79  + 459 : begin {REGofMAX1DataOut_F4_74[21:0] , REGofMAX1DataOut_F4_75[33:24] } <= AXIinput ; end 
80  + 459 : begin {REGofMAX1DataOut_F4_75[23:0] , REGofMAX1DataOut_F4_76[33:26] } <= AXIinput ; end 
81  + 459 : begin {REGofMAX1DataOut_F4_76[25:0] , REGofMAX1DataOut_F4_77[33:28] } <= AXIinput ; end 
82  + 459 : begin {REGofMAX1DataOut_F4_77[27:0] , REGofMAX1DataOut_F4_78[33:30] } <= AXIinput ; end 
83  + 459 : begin {REGofMAX1DataOut_F4_78[29:0] , REGofMAX1DataOut_F4_79[33:32] } <= AXIinput ; end 
84  + 459 : begin {REGofMAX1DataOut_F4_79[31:0] } <= AXIinput ; end 
85  + 459 : begin {REGofMAX1DataOut_F4_80[33:2] } <= AXIinput ; end 
86  + 459 : begin {REGofMAX1DataOut_F4_80[1:0], REGofMAX1DataOut_F4_81[33:4] } <= AXIinput ; end 
87  + 459 : begin {REGofMAX1DataOut_F4_81[3:0] , REGofMAX1DataOut_F4_82[33:6]  } <= AXIinput ; end 
88  + 459 : begin {REGofMAX1DataOut_F4_82[5:0] , REGofMAX1DataOut_F4_83[33:8]  } <= AXIinput ; end 
89  + 459 : begin {REGofMAX1DataOut_F4_83[7:0] , REGofMAX1DataOut_F4_84[33:10]  } <= AXIinput ; end 
90  + 459 : begin {REGofMAX1DataOut_F4_84[9:0] , REGofMAX1DataOut_F4_85[33:12]  } <= AXIinput ; end 
91  + 459 : begin {REGofMAX1DataOut_F4_85[11:0] , REGofMAX1DataOut_F4_86[33:14] } <= AXIinput ; end  
92  + 459 : begin {REGofMAX1DataOut_F4_86[13:0] , REGofMAX1DataOut_F4_87[33:16] } <= AXIinput ; end 
93  + 459 : begin {REGofMAX1DataOut_F4_87[15:0] , REGofMAX1DataOut_F4_88[33:18] } <= AXIinput ; end 
94  + 459 : begin {REGofMAX1DataOut_F4_88[17:0] , REGofMAX1DataOut_F4_89[33:20] } <= AXIinput ; end 
95  + 459 : begin {REGofMAX1DataOut_F4_89[19:0] , REGofMAX1DataOut_F4_90[33:22] } <= AXIinput ; end 
96  + 459 : begin {REGofMAX1DataOut_F4_90[21:0] , REGofMAX1DataOut_F4_91[33:24] } <= AXIinput ; end 
97  + 459 : begin {REGofMAX1DataOut_F4_91[23:0] , REGofMAX1DataOut_F4_92[33:26] } <= AXIinput ; end 
98  + 459 : begin {REGofMAX1DataOut_F4_92[25:0] , REGofMAX1DataOut_F4_93[33:28] } <= AXIinput ; end 
99  + 459 : begin {REGofMAX1DataOut_F4_93[27:0] , REGofMAX1DataOut_F4_94[33:30] } <= AXIinput ; end 
100  + 459 : begin {REGofMAX1DataOut_F4_94[29:0] , REGofMAX1DataOut_F4_95[33:32] } <= AXIinput ; end 
101  + 459 : begin {REGofMAX1DataOut_F4_95[31:0] } <= AXIinput ; end 
102  + 459 : begin {REGofMAX1DataOut_F4_96[33:2] } <= AXIinput ; end 
103  + 459 : begin {REGofMAX1DataOut_F4_96[1:0], REGofMAX1DataOut_F4_97[33:4] } <= AXIinput ; end 
104  + 459 : begin {REGofMAX1DataOut_F4_97[3:0] , REGofMAX1DataOut_F4_98[33:6]  } <= AXIinput ; end 
105  + 459 : begin {REGofMAX1DataOut_F4_98[5:0] , REGofMAX1DataOut_F4_99[33:8]  } <= AXIinput ; end  
106  + 459 : begin {REGofMAX1DataOut_F4_99[7:0] , REGofMAX1DataOut_F4_100[33:10]  } <= AXIinput ; end 
107  + 459 : begin {REGofMAX1DataOut_F4_100[9:0] , REGofMAX1DataOut_F4_101[33:12]  } <= AXIinput ; end 
108  + 459 : begin {REGofMAX1DataOut_F4_101[11:0] , REGofMAX1DataOut_F4_102[33:14] } <= AXIinput ; end  
109  + 459 : begin {REGofMAX1DataOut_F4_102[13:0] , REGofMAX1DataOut_F4_103[33:16] } <= AXIinput ; end 
110  + 459 : begin {REGofMAX1DataOut_F4_103[15:0] , REGofMAX1DataOut_F4_104[33:18] } <= AXIinput ; end 
111  + 459 : begin {REGofMAX1DataOut_F4_104[17:0] , REGofMAX1DataOut_F4_105[33:20] } <= AXIinput ; end 
112  + 459 : begin {REGofMAX1DataOut_F4_105[19:0] , REGofMAX1DataOut_F4_106[33:22] } <= AXIinput ; end 
113  + 459 : begin {REGofMAX1DataOut_F4_106[21:0] , REGofMAX1DataOut_F4_107[33:24] } <= AXIinput ; end 
114  + 459 : begin {REGofMAX1DataOut_F4_107[23:0] , REGofMAX1DataOut_F4_108[33:26] } <= AXIinput ; end 
115  + 459 : begin {REGofMAX1DataOut_F4_108[25:0] , REGofMAX1DataOut_F4_109[33:28] } <= AXIinput ; end 
116  + 459 : begin {REGofMAX1DataOut_F4_109[27:0] , REGofMAX1DataOut_F4_110[33:30] } <= AXIinput ; end 
117  + 459 : begin {REGofMAX1DataOut_F4_110[29:0] , REGofMAX1DataOut_F4_111[33:32] } <= AXIinput ; end 
118  + 459 : begin {REGofMAX1DataOut_F4_111[31:0] } <= AXIinput ; end 
119  + 459 : begin {REGofMAX1DataOut_F4_112[33:2] } <= AXIinput ; end 
120  + 459 : begin {REGofMAX1DataOut_F4_112[1:0], REGofMAX1DataOut_F4_113[33:4] } <= AXIinput ; end 
121  + 459 : begin {REGofMAX1DataOut_F4_113[3:0] , REGofMAX1DataOut_F4_114[33:6]  } <= AXIinput ; end 
122  + 459 : begin {REGofMAX1DataOut_F4_114[5:0] , REGofMAX1DataOut_F4_115[33:8]  } <= AXIinput ; end 
123  + 459 : begin {REGofMAX1DataOut_F4_115[7:0] , REGofMAX1DataOut_F4_116[33:10]  } <= AXIinput ; end 
124  + 459 : begin {REGofMAX1DataOut_F4_116[9:0] , REGofMAX1DataOut_F4_117[33:12]  } <= AXIinput ; end 
125  + 459 : begin {REGofMAX1DataOut_F4_117[11:0] , REGofMAX1DataOut_F4_118[33:14] } <= AXIinput ; end 
126  + 459 : begin {REGofMAX1DataOut_F4_118[13:0] , REGofMAX1DataOut_F4_119[33:16] } <= AXIinput ; end 
127  + 459 : begin {REGofMAX1DataOut_F4_119[15:0] , REGofMAX1DataOut_F4_120[33:18] } <= AXIinput ; end 
128  + 459 : begin {REGofMAX1DataOut_F4_120[17:0] , REGofMAX1DataOut_F4_121[33:20] } <= AXIinput ; end 
129  + 459 : begin {REGofMAX1DataOut_F4_121[19:0] , REGofMAX1DataOut_F4_122[33:22] } <= AXIinput ; end 
130  + 459 : begin {REGofMAX1DataOut_F4_122[21:0] , REGofMAX1DataOut_F4_123[33:24] } <= AXIinput ; end 
131  + 459 : begin {REGofMAX1DataOut_F4_123[23:0] , REGofMAX1DataOut_F4_124[33:26] } <= AXIinput ; end 
132  + 459 : begin {REGofMAX1DataOut_F4_124[25:0] , REGofMAX1DataOut_F4_125[33:28] } <= AXIinput ; end 
133  + 459 : begin {REGofMAX1DataOut_F4_125[27:0] , REGofMAX1DataOut_F4_126[33:30] } <= AXIinput ; end 
134  + 459 : begin {REGofMAX1DataOut_F4_126[29:0] , REGofMAX1DataOut_F4_127[33:32] } <= AXIinput ; end 
135  + 459 : begin {REGofMAX1DataOut_F4_127[31:0] } <= AXIinput ; end 
136  + 459 : begin {REGofMAX1DataOut_F4_128[33:2] } <= AXIinput ; end 
137  + 459 : begin {REGofMAX1DataOut_F4_128[1:0], REGofMAX1DataOut_F4_129[33:4] } <= AXIinput ; end 
138  + 459 : begin {REGofMAX1DataOut_F4_129[3:0] , REGofMAX1DataOut_F4_130[33:6]  } <= AXIinput ; end 
139  + 459 : begin {REGofMAX1DataOut_F4_130[5:0] , REGofMAX1DataOut_F4_131[33:8]  } <= AXIinput ; end 
140  + 459 : begin {REGofMAX1DataOut_F4_131[7:0] , REGofMAX1DataOut_F4_132[33:10]  } <= AXIinput ; end 
141  + 459 : begin {REGofMAX1DataOut_F4_132[9:0] , REGofMAX1DataOut_F4_133[33:12]  } <= AXIinput ; end 
142  + 459 : begin {REGofMAX1DataOut_F4_133[11:0] , REGofMAX1DataOut_F4_134[33:14] } <= AXIinput ; end 
143  + 459 : begin {REGofMAX1DataOut_F4_134[13:0] , REGofMAX1DataOut_F4_135[33:16] } <= AXIinput ; end 
144  + 459 : begin {REGofMAX1DataOut_F4_135[15:0] , REGofMAX1DataOut_F4_136[33:18] } <= AXIinput ; end 
145  + 459 : begin {REGofMAX1DataOut_F4_136[17:0] , REGofMAX1DataOut_F4_137[33:20] } <= AXIinput ; end 
146  + 459 : begin {REGofMAX1DataOut_F4_137[19:0] , REGofMAX1DataOut_F4_138[33:22] } <= AXIinput ; end 
147  + 459 : begin {REGofMAX1DataOut_F4_138[21:0] , REGofMAX1DataOut_F4_139[33:24] } <= AXIinput ; end 
148  + 459 : begin {REGofMAX1DataOut_F4_139[23:0] , REGofMAX1DataOut_F4_140[33:26] } <= AXIinput ; end 
149  + 459 : begin {REGofMAX1DataOut_F4_140[25:0] , REGofMAX1DataOut_F4_141[33:28] } <= AXIinput ; end 
150  + 459 : begin {REGofMAX1DataOut_F4_141[27:0] , REGofMAX1DataOut_F4_142[33:30] } <= AXIinput ; end 
151  + 459 : begin {REGofMAX1DataOut_F4_142[29:0] , REGofMAX1DataOut_F4_143[33:32] } <= AXIinput ; end 
152  + 459 : begin {REGofMAX1DataOut_F4_143[31:0] } <= AXIinput ; end 

612  : begin L0FINISH<= 1; end 
default: begin L0FINISH<= 1; end 
endcase


end
end

endmodule


//module happy(clk, rst_Controller,  AXIinput, AXIoutput, inputAXIstart  );
//input clk, rst_Controller, inputAXIstart;

module happy(clk,  AXIinput, AXIoutput  );
input clk;
input [31:0] AXIinput;
output [31:0] AXIoutput;
wire inputAXIstart;
assign inputAXIstart = 1'b1;
reg helpme = 1'b0;
always @(posedge clk) begin
helpme =  (inputAXIstart)? 1'b1:0;
end

//wire Conv2LayerStart;
wire MAX2LayerFinish;


//main_fsm_3_scenario31 MAINCONTROLLER_third_integration(clk, rst_Controller , MAX2LayerFinish, Conv2LayerStart);


wire [33:0]  REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143; 
wire [33:0]  REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143; 
wire [33:0]  REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143; 
wire [33:0]  REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143; 

wire [33:0] MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 ;

//wire L0FINISH; 
wire Conv2LayerStart;

AXIinputFromARM_3_1 axiINmodule (clk, AXIinput, helpme , Conv2LayerStart,
REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143 
);

MERGEHOPE_L3_L4  HOPE_3_4 (clk, Conv2LayerStart, MAX2LayerFinish
,REGofMAX1DataOut_F1_0,REGofMAX1DataOut_F1_1,REGofMAX1DataOut_F1_2,REGofMAX1DataOut_F1_3,REGofMAX1DataOut_F1_4,REGofMAX1DataOut_F1_5,REGofMAX1DataOut_F1_6,REGofMAX1DataOut_F1_7,REGofMAX1DataOut_F1_8,REGofMAX1DataOut_F1_9,REGofMAX1DataOut_F1_10,REGofMAX1DataOut_F1_11,REGofMAX1DataOut_F1_12,REGofMAX1DataOut_F1_13,REGofMAX1DataOut_F1_14,REGofMAX1DataOut_F1_15,REGofMAX1DataOut_F1_16,REGofMAX1DataOut_F1_17,REGofMAX1DataOut_F1_18,REGofMAX1DataOut_F1_19,REGofMAX1DataOut_F1_20,REGofMAX1DataOut_F1_21,REGofMAX1DataOut_F1_22,REGofMAX1DataOut_F1_23,REGofMAX1DataOut_F1_24,REGofMAX1DataOut_F1_25,REGofMAX1DataOut_F1_26,REGofMAX1DataOut_F1_27,REGofMAX1DataOut_F1_28,REGofMAX1DataOut_F1_29,REGofMAX1DataOut_F1_30,REGofMAX1DataOut_F1_31,REGofMAX1DataOut_F1_32,REGofMAX1DataOut_F1_33,REGofMAX1DataOut_F1_34,REGofMAX1DataOut_F1_35,REGofMAX1DataOut_F1_36,REGofMAX1DataOut_F1_37,REGofMAX1DataOut_F1_38,REGofMAX1DataOut_F1_39,REGofMAX1DataOut_F1_40,REGofMAX1DataOut_F1_41,REGofMAX1DataOut_F1_42,REGofMAX1DataOut_F1_43,REGofMAX1DataOut_F1_44,REGofMAX1DataOut_F1_45,REGofMAX1DataOut_F1_46,REGofMAX1DataOut_F1_47,REGofMAX1DataOut_F1_48,REGofMAX1DataOut_F1_49,REGofMAX1DataOut_F1_50,REGofMAX1DataOut_F1_51,REGofMAX1DataOut_F1_52,REGofMAX1DataOut_F1_53,REGofMAX1DataOut_F1_54,REGofMAX1DataOut_F1_55,REGofMAX1DataOut_F1_56,REGofMAX1DataOut_F1_57,REGofMAX1DataOut_F1_58,REGofMAX1DataOut_F1_59,REGofMAX1DataOut_F1_60,REGofMAX1DataOut_F1_61,REGofMAX1DataOut_F1_62,REGofMAX1DataOut_F1_63,REGofMAX1DataOut_F1_64,REGofMAX1DataOut_F1_65,REGofMAX1DataOut_F1_66,REGofMAX1DataOut_F1_67,REGofMAX1DataOut_F1_68,REGofMAX1DataOut_F1_69,REGofMAX1DataOut_F1_70,REGofMAX1DataOut_F1_71,REGofMAX1DataOut_F1_72,REGofMAX1DataOut_F1_73,REGofMAX1DataOut_F1_74,REGofMAX1DataOut_F1_75,REGofMAX1DataOut_F1_76,REGofMAX1DataOut_F1_77,REGofMAX1DataOut_F1_78,REGofMAX1DataOut_F1_79,REGofMAX1DataOut_F1_80,REGofMAX1DataOut_F1_81,REGofMAX1DataOut_F1_82,REGofMAX1DataOut_F1_83,REGofMAX1DataOut_F1_84,REGofMAX1DataOut_F1_85,REGofMAX1DataOut_F1_86,REGofMAX1DataOut_F1_87,REGofMAX1DataOut_F1_88,REGofMAX1DataOut_F1_89,REGofMAX1DataOut_F1_90,REGofMAX1DataOut_F1_91,REGofMAX1DataOut_F1_92,REGofMAX1DataOut_F1_93,REGofMAX1DataOut_F1_94,REGofMAX1DataOut_F1_95,REGofMAX1DataOut_F1_96,REGofMAX1DataOut_F1_97,REGofMAX1DataOut_F1_98,REGofMAX1DataOut_F1_99,REGofMAX1DataOut_F1_100,REGofMAX1DataOut_F1_101,REGofMAX1DataOut_F1_102,REGofMAX1DataOut_F1_103,REGofMAX1DataOut_F1_104,REGofMAX1DataOut_F1_105,REGofMAX1DataOut_F1_106,REGofMAX1DataOut_F1_107,REGofMAX1DataOut_F1_108,REGofMAX1DataOut_F1_109,REGofMAX1DataOut_F1_110,REGofMAX1DataOut_F1_111,REGofMAX1DataOut_F1_112,REGofMAX1DataOut_F1_113,REGofMAX1DataOut_F1_114,REGofMAX1DataOut_F1_115,REGofMAX1DataOut_F1_116,REGofMAX1DataOut_F1_117,REGofMAX1DataOut_F1_118,REGofMAX1DataOut_F1_119,REGofMAX1DataOut_F1_120,REGofMAX1DataOut_F1_121,REGofMAX1DataOut_F1_122,REGofMAX1DataOut_F1_123,REGofMAX1DataOut_F1_124,REGofMAX1DataOut_F1_125,REGofMAX1DataOut_F1_126,REGofMAX1DataOut_F1_127,REGofMAX1DataOut_F1_128,REGofMAX1DataOut_F1_129,REGofMAX1DataOut_F1_130,REGofMAX1DataOut_F1_131,REGofMAX1DataOut_F1_132,REGofMAX1DataOut_F1_133,REGofMAX1DataOut_F1_134,REGofMAX1DataOut_F1_135,REGofMAX1DataOut_F1_136,REGofMAX1DataOut_F1_137,REGofMAX1DataOut_F1_138,REGofMAX1DataOut_F1_139,REGofMAX1DataOut_F1_140,REGofMAX1DataOut_F1_141,REGofMAX1DataOut_F1_142,REGofMAX1DataOut_F1_143
,REGofMAX1DataOut_F2_0,REGofMAX1DataOut_F2_1,REGofMAX1DataOut_F2_2,REGofMAX1DataOut_F2_3,REGofMAX1DataOut_F2_4,REGofMAX1DataOut_F2_5,REGofMAX1DataOut_F2_6,REGofMAX1DataOut_F2_7,REGofMAX1DataOut_F2_8,REGofMAX1DataOut_F2_9,REGofMAX1DataOut_F2_10,REGofMAX1DataOut_F2_11,REGofMAX1DataOut_F2_12,REGofMAX1DataOut_F2_13,REGofMAX1DataOut_F2_14,REGofMAX1DataOut_F2_15,REGofMAX1DataOut_F2_16,REGofMAX1DataOut_F2_17,REGofMAX1DataOut_F2_18,REGofMAX1DataOut_F2_19,REGofMAX1DataOut_F2_20,REGofMAX1DataOut_F2_21,REGofMAX1DataOut_F2_22,REGofMAX1DataOut_F2_23,REGofMAX1DataOut_F2_24,REGofMAX1DataOut_F2_25,REGofMAX1DataOut_F2_26,REGofMAX1DataOut_F2_27,REGofMAX1DataOut_F2_28,REGofMAX1DataOut_F2_29,REGofMAX1DataOut_F2_30,REGofMAX1DataOut_F2_31,REGofMAX1DataOut_F2_32,REGofMAX1DataOut_F2_33,REGofMAX1DataOut_F2_34,REGofMAX1DataOut_F2_35,REGofMAX1DataOut_F2_36,REGofMAX1DataOut_F2_37,REGofMAX1DataOut_F2_38,REGofMAX1DataOut_F2_39,REGofMAX1DataOut_F2_40,REGofMAX1DataOut_F2_41,REGofMAX1DataOut_F2_42,REGofMAX1DataOut_F2_43,REGofMAX1DataOut_F2_44,REGofMAX1DataOut_F2_45,REGofMAX1DataOut_F2_46,REGofMAX1DataOut_F2_47,REGofMAX1DataOut_F2_48,REGofMAX1DataOut_F2_49,REGofMAX1DataOut_F2_50,REGofMAX1DataOut_F2_51,REGofMAX1DataOut_F2_52,REGofMAX1DataOut_F2_53,REGofMAX1DataOut_F2_54,REGofMAX1DataOut_F2_55,REGofMAX1DataOut_F2_56,REGofMAX1DataOut_F2_57,REGofMAX1DataOut_F2_58,REGofMAX1DataOut_F2_59,REGofMAX1DataOut_F2_60,REGofMAX1DataOut_F2_61,REGofMAX1DataOut_F2_62,REGofMAX1DataOut_F2_63,REGofMAX1DataOut_F2_64,REGofMAX1DataOut_F2_65,REGofMAX1DataOut_F2_66,REGofMAX1DataOut_F2_67,REGofMAX1DataOut_F2_68,REGofMAX1DataOut_F2_69,REGofMAX1DataOut_F2_70,REGofMAX1DataOut_F2_71,REGofMAX1DataOut_F2_72,REGofMAX1DataOut_F2_73,REGofMAX1DataOut_F2_74,REGofMAX1DataOut_F2_75,REGofMAX1DataOut_F2_76,REGofMAX1DataOut_F2_77,REGofMAX1DataOut_F2_78,REGofMAX1DataOut_F2_79,REGofMAX1DataOut_F2_80,REGofMAX1DataOut_F2_81,REGofMAX1DataOut_F2_82,REGofMAX1DataOut_F2_83,REGofMAX1DataOut_F2_84,REGofMAX1DataOut_F2_85,REGofMAX1DataOut_F2_86,REGofMAX1DataOut_F2_87,REGofMAX1DataOut_F2_88,REGofMAX1DataOut_F2_89,REGofMAX1DataOut_F2_90,REGofMAX1DataOut_F2_91,REGofMAX1DataOut_F2_92,REGofMAX1DataOut_F2_93,REGofMAX1DataOut_F2_94,REGofMAX1DataOut_F2_95,REGofMAX1DataOut_F2_96,REGofMAX1DataOut_F2_97,REGofMAX1DataOut_F2_98,REGofMAX1DataOut_F2_99,REGofMAX1DataOut_F2_100,REGofMAX1DataOut_F2_101,REGofMAX1DataOut_F2_102,REGofMAX1DataOut_F2_103,REGofMAX1DataOut_F2_104,REGofMAX1DataOut_F2_105,REGofMAX1DataOut_F2_106,REGofMAX1DataOut_F2_107,REGofMAX1DataOut_F2_108,REGofMAX1DataOut_F2_109,REGofMAX1DataOut_F2_110,REGofMAX1DataOut_F2_111,REGofMAX1DataOut_F2_112,REGofMAX1DataOut_F2_113,REGofMAX1DataOut_F2_114,REGofMAX1DataOut_F2_115,REGofMAX1DataOut_F2_116,REGofMAX1DataOut_F2_117,REGofMAX1DataOut_F2_118,REGofMAX1DataOut_F2_119,REGofMAX1DataOut_F2_120,REGofMAX1DataOut_F2_121,REGofMAX1DataOut_F2_122,REGofMAX1DataOut_F2_123,REGofMAX1DataOut_F2_124,REGofMAX1DataOut_F2_125,REGofMAX1DataOut_F2_126,REGofMAX1DataOut_F2_127,REGofMAX1DataOut_F2_128,REGofMAX1DataOut_F2_129,REGofMAX1DataOut_F2_130,REGofMAX1DataOut_F2_131,REGofMAX1DataOut_F2_132,REGofMAX1DataOut_F2_133,REGofMAX1DataOut_F2_134,REGofMAX1DataOut_F2_135,REGofMAX1DataOut_F2_136,REGofMAX1DataOut_F2_137,REGofMAX1DataOut_F2_138,REGofMAX1DataOut_F2_139,REGofMAX1DataOut_F2_140,REGofMAX1DataOut_F2_141,REGofMAX1DataOut_F2_142,REGofMAX1DataOut_F2_143 
,REGofMAX1DataOut_F3_0,REGofMAX1DataOut_F3_1,REGofMAX1DataOut_F3_2,REGofMAX1DataOut_F3_3,REGofMAX1DataOut_F3_4,REGofMAX1DataOut_F3_5,REGofMAX1DataOut_F3_6,REGofMAX1DataOut_F3_7,REGofMAX1DataOut_F3_8,REGofMAX1DataOut_F3_9,REGofMAX1DataOut_F3_10,REGofMAX1DataOut_F3_11,REGofMAX1DataOut_F3_12,REGofMAX1DataOut_F3_13,REGofMAX1DataOut_F3_14,REGofMAX1DataOut_F3_15,REGofMAX1DataOut_F3_16,REGofMAX1DataOut_F3_17,REGofMAX1DataOut_F3_18,REGofMAX1DataOut_F3_19,REGofMAX1DataOut_F3_20,REGofMAX1DataOut_F3_21,REGofMAX1DataOut_F3_22,REGofMAX1DataOut_F3_23,REGofMAX1DataOut_F3_24,REGofMAX1DataOut_F3_25,REGofMAX1DataOut_F3_26,REGofMAX1DataOut_F3_27,REGofMAX1DataOut_F3_28,REGofMAX1DataOut_F3_29,REGofMAX1DataOut_F3_30,REGofMAX1DataOut_F3_31,REGofMAX1DataOut_F3_32,REGofMAX1DataOut_F3_33,REGofMAX1DataOut_F3_34,REGofMAX1DataOut_F3_35,REGofMAX1DataOut_F3_36,REGofMAX1DataOut_F3_37,REGofMAX1DataOut_F3_38,REGofMAX1DataOut_F3_39,REGofMAX1DataOut_F3_40,REGofMAX1DataOut_F3_41,REGofMAX1DataOut_F3_42,REGofMAX1DataOut_F3_43,REGofMAX1DataOut_F3_44,REGofMAX1DataOut_F3_45,REGofMAX1DataOut_F3_46,REGofMAX1DataOut_F3_47,REGofMAX1DataOut_F3_48,REGofMAX1DataOut_F3_49,REGofMAX1DataOut_F3_50,REGofMAX1DataOut_F3_51,REGofMAX1DataOut_F3_52,REGofMAX1DataOut_F3_53,REGofMAX1DataOut_F3_54,REGofMAX1DataOut_F3_55,REGofMAX1DataOut_F3_56,REGofMAX1DataOut_F3_57,REGofMAX1DataOut_F3_58,REGofMAX1DataOut_F3_59,REGofMAX1DataOut_F3_60,REGofMAX1DataOut_F3_61,REGofMAX1DataOut_F3_62,REGofMAX1DataOut_F3_63,REGofMAX1DataOut_F3_64,REGofMAX1DataOut_F3_65,REGofMAX1DataOut_F3_66,REGofMAX1DataOut_F3_67,REGofMAX1DataOut_F3_68,REGofMAX1DataOut_F3_69,REGofMAX1DataOut_F3_70,REGofMAX1DataOut_F3_71,REGofMAX1DataOut_F3_72,REGofMAX1DataOut_F3_73,REGofMAX1DataOut_F3_74,REGofMAX1DataOut_F3_75,REGofMAX1DataOut_F3_76,REGofMAX1DataOut_F3_77,REGofMAX1DataOut_F3_78,REGofMAX1DataOut_F3_79,REGofMAX1DataOut_F3_80,REGofMAX1DataOut_F3_81,REGofMAX1DataOut_F3_82,REGofMAX1DataOut_F3_83,REGofMAX1DataOut_F3_84,REGofMAX1DataOut_F3_85,REGofMAX1DataOut_F3_86,REGofMAX1DataOut_F3_87,REGofMAX1DataOut_F3_88,REGofMAX1DataOut_F3_89,REGofMAX1DataOut_F3_90,REGofMAX1DataOut_F3_91,REGofMAX1DataOut_F3_92,REGofMAX1DataOut_F3_93,REGofMAX1DataOut_F3_94,REGofMAX1DataOut_F3_95,REGofMAX1DataOut_F3_96,REGofMAX1DataOut_F3_97,REGofMAX1DataOut_F3_98,REGofMAX1DataOut_F3_99,REGofMAX1DataOut_F3_100,REGofMAX1DataOut_F3_101,REGofMAX1DataOut_F3_102,REGofMAX1DataOut_F3_103,REGofMAX1DataOut_F3_104,REGofMAX1DataOut_F3_105,REGofMAX1DataOut_F3_106,REGofMAX1DataOut_F3_107,REGofMAX1DataOut_F3_108,REGofMAX1DataOut_F3_109,REGofMAX1DataOut_F3_110,REGofMAX1DataOut_F3_111,REGofMAX1DataOut_F3_112,REGofMAX1DataOut_F3_113,REGofMAX1DataOut_F3_114,REGofMAX1DataOut_F3_115,REGofMAX1DataOut_F3_116,REGofMAX1DataOut_F3_117,REGofMAX1DataOut_F3_118,REGofMAX1DataOut_F3_119,REGofMAX1DataOut_F3_120,REGofMAX1DataOut_F3_121,REGofMAX1DataOut_F3_122,REGofMAX1DataOut_F3_123,REGofMAX1DataOut_F3_124,REGofMAX1DataOut_F3_125,REGofMAX1DataOut_F3_126,REGofMAX1DataOut_F3_127,REGofMAX1DataOut_F3_128,REGofMAX1DataOut_F3_129,REGofMAX1DataOut_F3_130,REGofMAX1DataOut_F3_131,REGofMAX1DataOut_F3_132,REGofMAX1DataOut_F3_133,REGofMAX1DataOut_F3_134,REGofMAX1DataOut_F3_135,REGofMAX1DataOut_F3_136,REGofMAX1DataOut_F3_137,REGofMAX1DataOut_F3_138,REGofMAX1DataOut_F3_139,REGofMAX1DataOut_F3_140,REGofMAX1DataOut_F3_141,REGofMAX1DataOut_F3_142,REGofMAX1DataOut_F3_143 
,REGofMAX1DataOut_F4_0,REGofMAX1DataOut_F4_1,REGofMAX1DataOut_F4_2,REGofMAX1DataOut_F4_3,REGofMAX1DataOut_F4_4,REGofMAX1DataOut_F4_5,REGofMAX1DataOut_F4_6,REGofMAX1DataOut_F4_7,REGofMAX1DataOut_F4_8,REGofMAX1DataOut_F4_9,REGofMAX1DataOut_F4_10,REGofMAX1DataOut_F4_11,REGofMAX1DataOut_F4_12,REGofMAX1DataOut_F4_13,REGofMAX1DataOut_F4_14,REGofMAX1DataOut_F4_15,REGofMAX1DataOut_F4_16,REGofMAX1DataOut_F4_17,REGofMAX1DataOut_F4_18,REGofMAX1DataOut_F4_19,REGofMAX1DataOut_F4_20,REGofMAX1DataOut_F4_21,REGofMAX1DataOut_F4_22,REGofMAX1DataOut_F4_23,REGofMAX1DataOut_F4_24,REGofMAX1DataOut_F4_25,REGofMAX1DataOut_F4_26,REGofMAX1DataOut_F4_27,REGofMAX1DataOut_F4_28,REGofMAX1DataOut_F4_29,REGofMAX1DataOut_F4_30,REGofMAX1DataOut_F4_31,REGofMAX1DataOut_F4_32,REGofMAX1DataOut_F4_33,REGofMAX1DataOut_F4_34,REGofMAX1DataOut_F4_35,REGofMAX1DataOut_F4_36,REGofMAX1DataOut_F4_37,REGofMAX1DataOut_F4_38,REGofMAX1DataOut_F4_39,REGofMAX1DataOut_F4_40,REGofMAX1DataOut_F4_41,REGofMAX1DataOut_F4_42,REGofMAX1DataOut_F4_43,REGofMAX1DataOut_F4_44,REGofMAX1DataOut_F4_45,REGofMAX1DataOut_F4_46,REGofMAX1DataOut_F4_47,REGofMAX1DataOut_F4_48,REGofMAX1DataOut_F4_49,REGofMAX1DataOut_F4_50,REGofMAX1DataOut_F4_51,REGofMAX1DataOut_F4_52,REGofMAX1DataOut_F4_53,REGofMAX1DataOut_F4_54,REGofMAX1DataOut_F4_55,REGofMAX1DataOut_F4_56,REGofMAX1DataOut_F4_57,REGofMAX1DataOut_F4_58,REGofMAX1DataOut_F4_59,REGofMAX1DataOut_F4_60,REGofMAX1DataOut_F4_61,REGofMAX1DataOut_F4_62,REGofMAX1DataOut_F4_63,REGofMAX1DataOut_F4_64,REGofMAX1DataOut_F4_65,REGofMAX1DataOut_F4_66,REGofMAX1DataOut_F4_67,REGofMAX1DataOut_F4_68,REGofMAX1DataOut_F4_69,REGofMAX1DataOut_F4_70,REGofMAX1DataOut_F4_71,REGofMAX1DataOut_F4_72,REGofMAX1DataOut_F4_73,REGofMAX1DataOut_F4_74,REGofMAX1DataOut_F4_75,REGofMAX1DataOut_F4_76,REGofMAX1DataOut_F4_77,REGofMAX1DataOut_F4_78,REGofMAX1DataOut_F4_79,REGofMAX1DataOut_F4_80,REGofMAX1DataOut_F4_81,REGofMAX1DataOut_F4_82,REGofMAX1DataOut_F4_83,REGofMAX1DataOut_F4_84,REGofMAX1DataOut_F4_85,REGofMAX1DataOut_F4_86,REGofMAX1DataOut_F4_87,REGofMAX1DataOut_F4_88,REGofMAX1DataOut_F4_89,REGofMAX1DataOut_F4_90,REGofMAX1DataOut_F4_91,REGofMAX1DataOut_F4_92,REGofMAX1DataOut_F4_93,REGofMAX1DataOut_F4_94,REGofMAX1DataOut_F4_95,REGofMAX1DataOut_F4_96,REGofMAX1DataOut_F4_97,REGofMAX1DataOut_F4_98,REGofMAX1DataOut_F4_99,REGofMAX1DataOut_F4_100,REGofMAX1DataOut_F4_101,REGofMAX1DataOut_F4_102,REGofMAX1DataOut_F4_103,REGofMAX1DataOut_F4_104,REGofMAX1DataOut_F4_105,REGofMAX1DataOut_F4_106,REGofMAX1DataOut_F4_107,REGofMAX1DataOut_F4_108,REGofMAX1DataOut_F4_109,REGofMAX1DataOut_F4_110,REGofMAX1DataOut_F4_111,REGofMAX1DataOut_F4_112,REGofMAX1DataOut_F4_113,REGofMAX1DataOut_F4_114,REGofMAX1DataOut_F4_115,REGofMAX1DataOut_F4_116,REGofMAX1DataOut_F4_117,REGofMAX1DataOut_F4_118,REGofMAX1DataOut_F4_119,REGofMAX1DataOut_F4_120,REGofMAX1DataOut_F4_121,REGofMAX1DataOut_F4_122,REGofMAX1DataOut_F4_123,REGofMAX1DataOut_F4_124,REGofMAX1DataOut_F4_125,REGofMAX1DataOut_F4_126,REGofMAX1DataOut_F4_127,REGofMAX1DataOut_F4_128,REGofMAX1DataOut_F4_129,REGofMAX1DataOut_F4_130,REGofMAX1DataOut_F4_131,REGofMAX1DataOut_F4_132,REGofMAX1DataOut_F4_133,REGofMAX1DataOut_F4_134,REGofMAX1DataOut_F4_135,REGofMAX1DataOut_F4_136,REGofMAX1DataOut_F4_137,REGofMAX1DataOut_F4_138,REGofMAX1DataOut_F4_139,REGofMAX1DataOut_F4_140,REGofMAX1DataOut_F4_141,REGofMAX1DataOut_F4_142,REGofMAX1DataOut_F4_143 
,MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 
 );
 
//reg outputstart ;
//always @(posedge clk) begin outputstart <= 1'b1; end
 
AXIoutputToARM_3_1 axiOUTmodule (clk, AXIoutput, MAX2LayerFinish , 
MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 
);

endmodule


module AXIoutputToARM_3_1 (clk, AXIoutput, outputAXIstart , 
MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 
);

input clk ,  outputAXIstart ;
output reg [31:0] AXIoutput;
input [33:0] MAX2Data2_OutF4_0,MAX2Data2_OutF4_1,MAX2Data2_OutF4_2,MAX2Data2_OutF4_3,MAX2Data2_OutF4_4,MAX2Data2_OutF4_5,MAX2Data2_OutF4_6,MAX2Data2_OutF4_7,MAX2Data2_OutF4_8,MAX2Data2_OutF4_9,MAX2Data2_OutF4_10,MAX2Data2_OutF4_11,MAX2Data2_OutF4_12,MAX2Data2_OutF4_13,MAX2Data2_OutF4_14,MAX2Data2_OutF4_15,MAX2Data2_OutF4_16,MAX2Data2_OutF4_17,MAX2Data2_OutF4_18,MAX2Data2_OutF4_19,MAX2Data2_OutF4_20,MAX2Data2_OutF4_21,MAX2Data2_OutF4_22,MAX2Data2_OutF4_23,MAX2Data2_OutF4_24 ;

reg L0FINISH;


wire [5:0] counter; 
COUNTER_LAYER_55_cycles TheCounter (clk, counter, outputAXIstart);
always @(posedge clk) 
begin 
if (outputAXIstart)
begin
case(counter)


0 : begin AXIoutput  <=  { MAX2Data2_OutF4_0[33:2]} ; end 
1 : begin AXIoutput  <=  { MAX2Data2_OutF4_0[1:0], MAX2Data2_OutF4_1[33:4]} ; end 
2 : begin AXIoutput  <=  { MAX2Data2_OutF4_1[3:0] , MAX2Data2_OutF4_2[33:6] } ; end 
3 : begin AXIoutput  <=  { MAX2Data2_OutF4_2[5:0] , MAX2Data2_OutF4_3[33:8] } ; end  
4 : begin AXIoutput  <=  { MAX2Data2_OutF4_3[7:0] , MAX2Data2_OutF4_4[33:10] } ; end 
5 : begin AXIoutput  <=  { MAX2Data2_OutF4_4[9:0] , MAX2Data2_OutF4_5[33:12] } ; end 
6 : begin AXIoutput  <=  { MAX2Data2_OutF4_5[11:0] , MAX2Data2_OutF4_6[33:14]} ; end 
7 : begin AXIoutput  <=  { MAX2Data2_OutF4_6[13:0] , MAX2Data2_OutF4_7[33:16]} ; end 
8 : begin AXIoutput  <=  { MAX2Data2_OutF4_7[15:0] , MAX2Data2_OutF4_8[33:18]} ; end 
9 : begin AXIoutput  <=  { MAX2Data2_OutF4_8[17:0] , MAX2Data2_OutF4_9[33:20]} ; end 
10 : begin AXIoutput  <=  { MAX2Data2_OutF4_9[19:0] , MAX2Data2_OutF4_10[33:22]} ; end 
11 : begin AXIoutput  <=  { MAX2Data2_OutF4_10[21:0] , MAX2Data2_OutF4_11[33:24]} ; end 
12 : begin AXIoutput  <=  { MAX2Data2_OutF4_11[23:0] , MAX2Data2_OutF4_12[33:26]} ; end 
13 : begin AXIoutput  <=  { MAX2Data2_OutF4_12[25:0] , MAX2Data2_OutF4_13[33:28]} ; end 
14 : begin AXIoutput  <=  { MAX2Data2_OutF4_13[27:0] , MAX2Data2_OutF4_14[33:30]} ; end 
15 : begin AXIoutput  <=  { MAX2Data2_OutF4_14[29:0] , MAX2Data2_OutF4_15[33:32]} ; end 
16 : begin AXIoutput  <=  { MAX2Data2_OutF4_15[31:0]} ; end 


17 : begin AXIoutput  <=  { MAX2Data2_OutF4_16[33:2]} ; end 
18 : begin AXIoutput  <=  { MAX2Data2_OutF4_16[1:0], MAX2Data2_OutF4_17[33:4]} ; end 
19 : begin AXIoutput  <=  { MAX2Data2_OutF4_17[3:0] , MAX2Data2_OutF4_18[33:6] } ; end 
20 : begin AXIoutput  <=  { MAX2Data2_OutF4_18[5:0] , MAX2Data2_OutF4_19[33:8] } ; end 
21 : begin AXIoutput  <=  { MAX2Data2_OutF4_19[7:0] , MAX2Data2_OutF4_20[33:10] } ; end 
22 : begin AXIoutput  <=  { MAX2Data2_OutF4_20[9:0] , MAX2Data2_OutF4_21[33:12] } ; end 
23 : begin AXIoutput  <=  { MAX2Data2_OutF4_21[11:0] , MAX2Data2_OutF4_22[33:14]} ; end 
24 : begin AXIoutput  <=  { MAX2Data2_OutF4_22[13:0] , MAX2Data2_OutF4_23[33:16]} ; end 
25 : begin AXIoutput  <=  { MAX2Data2_OutF4_23[15:0] , MAX2Data2_OutF4_24[33:18]} ; end  
26 : begin AXIoutput  <=  { MAX2Data2_OutF4_24[17:0] , 14'bxxxxxxxxxxxxxx} ; end 


27  : begin L0FINISH<= 1; end 
default: begin L0FINISH<= 1; end 
endcase
end
end


endmodule



module COUNTER_LAYER_55_cycles (clk, count_temp, AXIstart);

input clk;
input AXIstart;
output reg [5:0] count_temp;
initial begin count_temp <=6'b000000; end
always @ (posedge clk)
begin 
if(AXIstart)
count_temp <= count_temp +6'b000001;
end

endmodule



module COUNTER_LAYER_1200_cycles (clk, count_temp, AXIstart);

input clk;
input AXIstart;
output reg [10:0] count_temp;
initial begin count_temp <=11'b00000000000; end
always @ (posedge clk)
begin 
if(AXIstart)
count_temp <= count_temp +11'b00000000001;
end

endmodule































